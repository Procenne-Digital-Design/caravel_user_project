VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1500.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 1496.000 2.210 1500.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1496.000 113.070 1500.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 1496.000 124.110 1500.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 1496.000 135.150 1500.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 1496.000 146.650 1500.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 1496.000 157.690 1500.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 1496.000 168.730 1500.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 1496.000 179.770 1500.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 1496.000 190.810 1500.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 1496.000 201.850 1500.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1496.000 212.890 1500.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 1496.000 13.250 1500.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 1496.000 224.390 1500.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1496.000 235.430 1500.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 1496.000 246.470 1500.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 1496.000 257.510 1500.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 1496.000 268.550 1500.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 1496.000 279.590 1500.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 1496.000 291.090 1500.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 1496.000 302.130 1500.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 1496.000 313.170 1500.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 1496.000 324.210 1500.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 1496.000 24.290 1500.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1496.000 335.250 1500.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 1496.000 346.290 1500.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 1496.000 357.330 1500.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 1496.000 368.830 1500.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 1496.000 379.870 1500.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 1496.000 390.910 1500.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 1496.000 401.950 1500.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 1496.000 412.990 1500.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 1496.000 35.330 1500.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 1496.000 46.370 1500.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 1496.000 57.410 1500.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 1496.000 68.450 1500.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 1496.000 79.950 1500.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 1496.000 90.990 1500.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 1496.000 102.030 1500.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 1496.000 5.890 1500.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 1496.000 116.750 1500.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 1496.000 127.790 1500.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1496.000 138.830 1500.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 1496.000 150.330 1500.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1496.000 161.370 1500.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 1496.000 172.410 1500.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 1496.000 183.450 1500.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 1496.000 194.490 1500.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 1496.000 205.530 1500.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 1496.000 217.030 1500.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 1496.000 16.930 1500.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 1496.000 228.070 1500.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 1496.000 239.110 1500.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 1496.000 250.150 1500.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1496.000 261.190 1500.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 1496.000 272.230 1500.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 1496.000 283.270 1500.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 1496.000 294.770 1500.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 1496.000 305.810 1500.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 1496.000 316.850 1500.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 1496.000 327.890 1500.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 1496.000 27.970 1500.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 1496.000 338.930 1500.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 1496.000 349.970 1500.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 1496.000 361.470 1500.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 1496.000 372.510 1500.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1496.000 383.550 1500.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 1496.000 394.590 1500.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 1496.000 405.630 1500.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 1496.000 416.670 1500.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1496.000 39.010 1500.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 1496.000 50.050 1500.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 1496.000 61.090 1500.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 1496.000 72.130 1500.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 1496.000 83.630 1500.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 1496.000 94.670 1500.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 1496.000 105.710 1500.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 1496.000 9.570 1500.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 1496.000 120.430 1500.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 1496.000 131.470 1500.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 1496.000 142.510 1500.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 1496.000 154.010 1500.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 1496.000 165.050 1500.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 1496.000 176.090 1500.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 1496.000 187.130 1500.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 1496.000 198.170 1500.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 1496.000 209.210 1500.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 1496.000 220.710 1500.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 1496.000 20.610 1500.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 1496.000 231.750 1500.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 1496.000 242.790 1500.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 1496.000 253.830 1500.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 1496.000 264.870 1500.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 1496.000 275.910 1500.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1496.000 286.950 1500.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 1496.000 298.450 1500.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1496.000 309.490 1500.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 1496.000 320.530 1500.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 1496.000 331.570 1500.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 1496.000 31.650 1500.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 1496.000 342.610 1500.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 1496.000 353.650 1500.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 1496.000 365.150 1500.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 1496.000 376.190 1500.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 1496.000 387.230 1500.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 1496.000 398.270 1500.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 1496.000 409.310 1500.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 1496.000 420.350 1500.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 1496.000 42.690 1500.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 1496.000 53.730 1500.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1496.000 64.770 1500.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 1496.000 76.270 1500.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1496.000 87.310 1500.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 1496.000 98.350 1500.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 1496.000 109.390 1500.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 4.800 1000.000 5.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1324.000 1000.000 1324.600 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1345.080 1000.000 1345.680 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 1496.000 898.290 1500.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1355.280 1000.000 1355.880 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 1496.000 909.330 1500.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1366.160 1000.000 1366.760 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 1496.000 920.370 1500.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 0.000 948.890 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 1496.000 516.950 1500.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 1496.000 931.870 1500.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 1496.000 939.230 1500.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 1496.000 946.590 1500.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1398.120 1000.000 1398.720 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.760 4.000 1414.360 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 1496.000 957.630 1500.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.160 4.000 1434.760 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1444.360 4.000 1444.960 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1440.960 1000.000 1441.560 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 323.720 1000.000 324.320 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1464.080 4.000 1464.680 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 0.000 973.270 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 1496.000 979.710 1500.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.280 4.000 1474.880 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1484.480 4.000 1485.080 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 1496.000 994.430 1500.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1494.000 1000.000 1494.600 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 1496.000 524.310 1500.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 1496.000 542.710 1500.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 472.640 1000.000 473.240 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 1496.000 576.290 1500.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 525.680 1000.000 526.280 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 557.640 1000.000 558.240 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 568.520 1000.000 569.120 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 1496.000 627.810 1500.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 621.560 1000.000 622.160 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 695.680 1000.000 696.280 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 781.360 1000.000 781.960 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 1496.000 453.930 1500.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 1496.000 668.750 1500.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.280 4.000 709.880 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 1496.000 687.150 1500.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 866.360 1000.000 866.960 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 887.440 1000.000 888.040 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 908.520 1000.000 909.120 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 1496.000 709.230 1500.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 1496.000 717.050 1500.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1496.000 728.090 1500.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 1496.000 468.650 1500.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 1496.000 731.770 1500.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1025.480 1000.000 1026.080 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1036.360 1000.000 1036.960 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 4.000 900.960 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 910.560 4.000 911.160 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 1496.000 750.170 1500.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 1496.000 757.530 1500.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 1496.000 772.250 1500.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1496.000 779.610 1500.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 1496.000 786.970 1500.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.000 4.000 1001.600 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1021.400 4.000 1022.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 1496.000 798.470 1500.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1061.520 4.000 1062.120 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 1496.000 805.830 1500.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.920 4.000 1082.520 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1174.400 1000.000 1175.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 1496.000 813.190 1500.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1196.160 1000.000 1196.760 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 1496.000 820.550 1500.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 1496.000 824.230 1500.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 1496.000 827.910 1500.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 206.760 1000.000 207.360 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1217.240 1000.000 1217.840 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.330 0.000 871.610 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 1496.000 842.630 1500.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.280 4.000 1202.880 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1212.480 4.000 1213.080 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1232.880 4.000 1233.480 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 1496.000 502.230 1500.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 1496.000 857.350 1500.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 1496.000 865.170 1500.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1270.280 1000.000 1270.880 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1281.160 1000.000 1281.760 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 1496.000 872.530 1500.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1323.320 4.000 1323.920 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 1496.000 883.570 1500.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1333.520 4.000 1334.120 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 1496.000 887.250 1500.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1334.200 1000.000 1334.800 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 1496.000 890.930 1500.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.720 4.000 1344.320 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.730 1496.000 913.010 1500.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1377.040 1000.000 1377.640 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.470 0.000 944.750 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 1496.000 924.050 1500.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 1496.000 935.550 1500.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 1496.000 950.270 1500.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 0.000 961.310 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1403.560 4.000 1404.160 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 1496.000 953.950 1500.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1409.000 1000.000 1409.600 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 1496.000 964.990 1500.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1430.080 1000.000 1430.680 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1451.160 1000.000 1451.760 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 1496.000 520.630 1500.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 1496.000 976.030 1500.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 1496.000 983.390 1500.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 1496.000 987.070 1500.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 1496.000 990.750 1500.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 1496.000 998.110 1500.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1494.680 4.000 1495.280 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 1496.000 527.990 1500.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 397.840 1000.000 398.440 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 419.600 1000.000 420.200 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 1496.000 546.390 1500.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1496.000 579.970 1500.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 1496.000 591.010 1500.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 1496.000 616.770 1500.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 706.560 1000.000 707.160 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 78.920 1000.000 79.520 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 1496.000 690.830 1500.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 1496.000 694.510 1500.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 1496.000 698.190 1500.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.920 4.000 810.520 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 898.320 1000.000 898.920 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 1496.000 457.610 1500.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 830.320 4.000 830.920 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 919.400 1000.000 920.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 940.480 1000.000 941.080 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 951.360 1000.000 951.960 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 962.240 1000.000 962.840 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 983.320 1000.000 983.920 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 1496.000 735.450 1500.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1015.280 1000.000 1015.880 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.160 4.000 890.760 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1047.240 1000.000 1047.840 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1496.000 753.850 1500.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1068.320 1000.000 1068.920 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 1496.000 761.210 1500.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 1496.000 775.930 1500.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1079.200 1000.000 1079.800 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.280 4.000 981.880 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.800 4.000 991.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1111.160 1000.000 1111.760 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.200 4.000 1011.800 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1031.600 4.000 1032.200 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.120 4.000 1041.720 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.720 4.000 1072.320 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1143.120 1000.000 1143.720 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1153.320 1000.000 1153.920 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 0.000 850.910 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 1496.000 831.590 1500.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 216.960 1000.000 217.560 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1206.360 1000.000 1206.960 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1228.120 1000.000 1228.720 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1249.200 1000.000 1249.800 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1260.080 1000.000 1260.680 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1182.560 4.000 1183.160 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 0.000 883.570 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1222.680 4.000 1223.280 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1496.000 853.670 1500.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 1496.000 861.490 1500.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1273.000 4.000 1273.600 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 1496.000 868.850 1500.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.920 4.000 1303.520 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1313.120 4.000 1313.720 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 1496.000 879.890 1500.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1302.240 1000.000 1302.840 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1313.120 1000.000 1313.720 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 15.000 1000.000 15.600 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 0.000 920.370 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 0.000 928.650 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 1496.000 894.610 1500.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 1496.000 901.970 1500.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 1496.000 905.650 1500.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 1496.000 916.690 1500.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1387.240 1000.000 1387.840 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1496.000 927.730 1500.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 312.840 1000.000 313.440 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 0.000 953.030 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 1496.000 942.910 1500.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 0.000 957.170 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1423.960 4.000 1424.560 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 1496.000 961.310 1500.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1419.200 1000.000 1419.800 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 1496.000 968.670 1500.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1453.880 4.000 1454.480 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 1496.000 972.350 1500.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1462.040 1000.000 1462.640 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1472.920 1000.000 1473.520 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 0.000 981.550 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 0.000 993.970 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1483.120 1000.000 1483.720 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 0.000 998.110 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 355.680 1000.000 356.280 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 1496.000 535.350 1500.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 451.560 1000.000 452.160 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 504.600 1000.000 505.200 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 1496.000 583.650 1500.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 1496.000 446.570 1500.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 1496.000 598.370 1500.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 1496.000 620.450 1500.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 589.600 1000.000 590.200 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 632.440 1000.000 633.040 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 717.440 1000.000 718.040 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 749.400 1000.000 750.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 1496.000 661.390 1500.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 759.600 4.000 760.200 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 4.000 780.600 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 876.560 1000.000 877.160 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 1496.000 701.870 1500.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 1496.000 705.550 1500.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 930.280 1000.000 930.880 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 1496.000 712.910 1500.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 0.000 761.210 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 972.440 1000.000 973.040 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 1496.000 720.730 1500.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 1496.000 724.410 1500.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 994.200 1000.000 994.800 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1004.400 1000.000 1005.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 121.760 1000.000 122.360 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 1496.000 739.130 1500.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 1496.000 742.810 1500.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 1496.000 746.490 1500.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1057.440 1000.000 1058.040 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 1496.000 764.890 1500.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 1496.000 768.570 1500.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 153.720 1000.000 154.320 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 940.480 4.000 941.080 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 1496.000 783.290 1500.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1089.400 1000.000 1090.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1100.280 1000.000 1100.880 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 1496.000 791.110 1500.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1121.360 1000.000 1121.960 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 1496.000 794.790 1500.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1051.320 4.000 1051.920 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1132.240 1000.000 1132.840 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1496.000 802.150 1500.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 1496.000 809.510 1500.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1164.200 1000.000 1164.800 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1185.280 1000.000 1185.880 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 1496.000 816.870 1500.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 227.840 1000.000 228.440 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 1496.000 835.270 1500.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 1496.000 838.950 1500.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1238.320 1000.000 1238.920 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1172.360 4.000 1172.960 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1192.760 4.000 1193.360 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 1496.000 846.310 1500.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 1496.000 849.990 1500.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1252.600 4.000 1253.200 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1262.800 4.000 1263.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1283.200 4.000 1283.800 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1292.040 1000.000 1292.640 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1496.000 876.210 1500.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 0.000 904.270 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 0.000 907.950 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END la_oenb[9]
  PIN sram_addr_a[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 1496.000 431.850 1500.000 ;
    END
  END sram_addr_a[0]
  PIN sram_addr_a[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 36.080 1000.000 36.680 ;
    END
  END sram_addr_a[1]
  PIN sram_addr_a[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END sram_addr_a[2]
  PIN sram_addr_a[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 1496.000 461.290 1500.000 ;
    END
  END sram_addr_a[3]
  PIN sram_addr_a[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 131.960 1000.000 132.560 ;
    END
  END sram_addr_a[4]
  PIN sram_addr_a[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END sram_addr_a[5]
  PIN sram_addr_a[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 174.800 1000.000 175.400 ;
    END
  END sram_addr_a[6]
  PIN sram_addr_a[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 238.720 1000.000 239.320 ;
    END
  END sram_addr_a[7]
  PIN sram_addr_a[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END sram_addr_a[8]
  PIN sram_addr_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END sram_addr_b[0]
  PIN sram_addr_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 46.960 1000.000 47.560 ;
    END
  END sram_addr_b[1]
  PIN sram_addr_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END sram_addr_b[2]
  PIN sram_addr_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 100.000 1000.000 100.600 ;
    END
  END sram_addr_b[3]
  PIN sram_addr_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END sram_addr_b[4]
  PIN sram_addr_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END sram_addr_b[5]
  PIN sram_addr_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 1496.000 490.730 1500.000 ;
    END
  END sram_addr_b[6]
  PIN sram_addr_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END sram_addr_b[7]
  PIN sram_addr_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 259.800 1000.000 260.400 ;
    END
  END sram_addr_b[8]
  PIN sram_csb_a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END sram_csb_a
  PIN sram_csb_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END sram_csb_b
  PIN sram_din_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END sram_din_b[0]
  PIN sram_din_b[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END sram_din_b[10]
  PIN sram_din_b[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END sram_din_b[11]
  PIN sram_din_b[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1496.000 531.670 1500.000 ;
    END
  END sram_din_b[12]
  PIN sram_din_b[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END sram_din_b[13]
  PIN sram_din_b[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 429.800 1000.000 430.400 ;
    END
  END sram_din_b[14]
  PIN sram_din_b[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END sram_din_b[15]
  PIN sram_din_b[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 1496.000 561.110 1500.000 ;
    END
  END sram_din_b[16]
  PIN sram_din_b[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 1496.000 568.470 1500.000 ;
    END
  END sram_din_b[17]
  PIN sram_din_b[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END sram_din_b[18]
  PIN sram_din_b[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END sram_din_b[19]
  PIN sram_din_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 57.840 1000.000 58.440 ;
    END
  END sram_din_b[1]
  PIN sram_din_b[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END sram_din_b[20]
  PIN sram_din_b[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 1496.000 605.730 1500.000 ;
    END
  END sram_din_b[21]
  PIN sram_din_b[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END sram_din_b[22]
  PIN sram_din_b[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 578.720 1000.000 579.320 ;
    END
  END sram_din_b[23]
  PIN sram_din_b[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 1496.000 638.850 1500.000 ;
    END
  END sram_din_b[24]
  PIN sram_din_b[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 642.640 1000.000 643.240 ;
    END
  END sram_din_b[25]
  PIN sram_din_b[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 674.600 1000.000 675.200 ;
    END
  END sram_din_b[26]
  PIN sram_din_b[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 727.640 1000.000 728.240 ;
    END
  END sram_din_b[27]
  PIN sram_din_b[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 1496.000 657.710 1500.000 ;
    END
  END sram_din_b[28]
  PIN sram_din_b[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 791.560 1000.000 792.160 ;
    END
  END sram_din_b[29]
  PIN sram_din_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END sram_din_b[2]
  PIN sram_din_b[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 1496.000 672.430 1500.000 ;
    END
  END sram_din_b[30]
  PIN sram_din_b[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 855.480 1000.000 856.080 ;
    END
  END sram_din_b[31]
  PIN sram_din_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END sram_din_b[3]
  PIN sram_din_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END sram_din_b[4]
  PIN sram_din_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END sram_din_b[5]
  PIN sram_din_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END sram_din_b[6]
  PIN sram_din_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END sram_din_b[7]
  PIN sram_din_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 1496.000 505.910 1500.000 ;
    END
  END sram_din_b[8]
  PIN sram_din_b[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 1496.000 513.270 1500.000 ;
    END
  END sram_din_b[9]
  PIN sram_dout_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 25.880 1000.000 26.480 ;
    END
  END sram_dout_a[0]
  PIN sram_dout_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END sram_dout_a[10]
  PIN sram_dout_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 334.600 1000.000 335.200 ;
    END
  END sram_dout_a[11]
  PIN sram_dout_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 365.880 1000.000 366.480 ;
    END
  END sram_dout_a[12]
  PIN sram_dout_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END sram_dout_a[13]
  PIN sram_dout_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END sram_dout_a[14]
  PIN sram_dout_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 1496.000 550.070 1500.000 ;
    END
  END sram_dout_a[15]
  PIN sram_dout_a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 1496.000 564.790 1500.000 ;
    END
  END sram_dout_a[16]
  PIN sram_dout_a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 1496.000 572.150 1500.000 ;
    END
  END sram_dout_a[17]
  PIN sram_dout_a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 1496.000 587.330 1500.000 ;
    END
  END sram_dout_a[18]
  PIN sram_dout_a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END sram_dout_a[19]
  PIN sram_dout_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 1496.000 450.250 1500.000 ;
    END
  END sram_dout_a[1]
  PIN sram_dout_a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 1496.000 602.050 1500.000 ;
    END
  END sram_dout_a[20]
  PIN sram_dout_a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END sram_dout_a[21]
  PIN sram_dout_a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 1496.000 624.130 1500.000 ;
    END
  END sram_dout_a[22]
  PIN sram_dout_a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END sram_dout_a[23]
  PIN sram_dout_a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 600.480 1000.000 601.080 ;
    END
  END sram_dout_a[24]
  PIN sram_dout_a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 653.520 1000.000 654.120 ;
    END
  END sram_dout_a[25]
  PIN sram_dout_a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 0.000 691.750 4.000 ;
    END
  END sram_dout_a[26]
  PIN sram_dout_a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1496.000 654.030 1500.000 ;
    END
  END sram_dout_a[27]
  PIN sram_dout_a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 0.000 708.310 4.000 ;
    END
  END sram_dout_a[28]
  PIN sram_dout_a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 802.440 1000.000 803.040 ;
    END
  END sram_dout_a[29]
  PIN sram_dout_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END sram_dout_a[2]
  PIN sram_dout_a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 834.400 1000.000 835.000 ;
    END
  END sram_dout_a[30]
  PIN sram_dout_a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 1496.000 683.470 1500.000 ;
    END
  END sram_dout_a[31]
  PIN sram_dout_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END sram_dout_a[3]
  PIN sram_dout_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 1496.000 472.330 1500.000 ;
    END
  END sram_dout_a[4]
  PIN sram_dout_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 1496.000 479.690 1500.000 ;
    END
  END sram_dout_a[5]
  PIN sram_dout_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 185.000 1000.000 185.600 ;
    END
  END sram_dout_a[6]
  PIN sram_dout_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END sram_dout_a[7]
  PIN sram_dout_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END sram_dout_a[8]
  PIN sram_dout_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 291.760 1000.000 292.360 ;
    END
  END sram_dout_a[9]
  PIN sram_mask_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 1496.000 435.530 1500.000 ;
    END
  END sram_mask_b[0]
  PIN sram_mask_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END sram_mask_b[1]
  PIN sram_mask_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END sram_mask_b[2]
  PIN sram_mask_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END sram_mask_b[3]
  PIN sram_web_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END sram_web_b
  PIN trng_buffer_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END trng_buffer_i[0]
  PIN trng_buffer_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END trng_buffer_i[10]
  PIN trng_buffer_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END trng_buffer_i[11]
  PIN trng_buffer_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END trng_buffer_i[12]
  PIN trng_buffer_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END trng_buffer_i[13]
  PIN trng_buffer_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 1496.000 539.030 1500.000 ;
    END
  END trng_buffer_i[14]
  PIN trng_buffer_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 1496.000 553.750 1500.000 ;
    END
  END trng_buffer_i[15]
  PIN trng_buffer_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 483.520 1000.000 484.120 ;
    END
  END trng_buffer_i[16]
  PIN trng_buffer_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END trng_buffer_i[17]
  PIN trng_buffer_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END trng_buffer_i[18]
  PIN trng_buffer_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 1496.000 594.690 1500.000 ;
    END
  END trng_buffer_i[19]
  PIN trng_buffer_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END trng_buffer_i[1]
  PIN trng_buffer_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 0.000 654.950 4.000 ;
    END
  END trng_buffer_i[20]
  PIN trng_buffer_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 1496.000 609.410 1500.000 ;
    END
  END trng_buffer_i[21]
  PIN trng_buffer_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END trng_buffer_i[22]
  PIN trng_buffer_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END trng_buffer_i[23]
  PIN trng_buffer_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END trng_buffer_i[24]
  PIN trng_buffer_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 664.400 1000.000 665.000 ;
    END
  END trng_buffer_i[25]
  PIN trng_buffer_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END trng_buffer_i[26]
  PIN trng_buffer_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END trng_buffer_i[27]
  PIN trng_buffer_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 759.600 1000.000 760.200 ;
    END
  END trng_buffer_i[28]
  PIN trng_buffer_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 813.320 1000.000 813.920 ;
    END
  END trng_buffer_i[29]
  PIN trng_buffer_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 89.800 1000.000 90.400 ;
    END
  END trng_buffer_i[2]
  PIN trng_buffer_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 844.600 1000.000 845.200 ;
    END
  END trng_buffer_i[30]
  PIN trng_buffer_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.200 4.000 739.800 ;
    END
  END trng_buffer_i[31]
  PIN trng_buffer_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END trng_buffer_i[3]
  PIN trng_buffer_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END trng_buffer_i[4]
  PIN trng_buffer_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 1496.000 483.370 1500.000 ;
    END
  END trng_buffer_i[5]
  PIN trng_buffer_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END trng_buffer_i[6]
  PIN trng_buffer_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END trng_buffer_i[7]
  PIN trng_buffer_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 270.680 1000.000 271.280 ;
    END
  END trng_buffer_i[8]
  PIN trng_buffer_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 302.640 1000.000 303.240 ;
    END
  END trng_buffer_i[9]
  PIN trng_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 1496.000 424.030 1500.000 ;
    END
  END trng_wb_ack_i
  PIN trng_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 1496.000 439.210 1500.000 ;
    END
  END trng_wb_adr_o[0]
  PIN trng_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 68.040 1000.000 68.640 ;
    END
  END trng_wb_adr_o[1]
  PIN trng_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END trng_wb_adr_o[2]
  PIN trng_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END trng_wb_adr_o[3]
  PIN trng_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 1496.000 476.010 1500.000 ;
    END
  END trng_wb_adr_o[4]
  PIN trng_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 163.920 1000.000 164.520 ;
    END
  END trng_wb_adr_o[5]
  PIN trng_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 1496.000 494.410 1500.000 ;
    END
  END trng_wb_adr_o[6]
  PIN trng_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END trng_wb_adr_o[7]
  PIN trng_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 280.880 1000.000 281.480 ;
    END
  END trng_wb_adr_o[8]
  PIN trng_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END trng_wb_cyc_o
  PIN trng_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END trng_wb_dat_i[0]
  PIN trng_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END trng_wb_dat_i[10]
  PIN trng_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 344.800 1000.000 345.400 ;
    END
  END trng_wb_dat_i[11]
  PIN trng_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 376.760 1000.000 377.360 ;
    END
  END trng_wb_dat_i[12]
  PIN trng_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END trng_wb_dat_i[13]
  PIN trng_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 440.680 1000.000 441.280 ;
    END
  END trng_wb_dat_i[14]
  PIN trng_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 461.760 1000.000 462.360 ;
    END
  END trng_wb_dat_i[15]
  PIN trng_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 493.720 1000.000 494.320 ;
    END
  END trng_wb_dat_i[16]
  PIN trng_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END trng_wb_dat_i[17]
  PIN trng_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END trng_wb_dat_i[18]
  PIN trng_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END trng_wb_dat_i[19]
  PIN trng_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END trng_wb_dat_i[1]
  PIN trng_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 536.560 1000.000 537.160 ;
    END
  END trng_wb_dat_i[20]
  PIN trng_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 1496.000 613.090 1500.000 ;
    END
  END trng_wb_dat_i[21]
  PIN trng_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END trng_wb_dat_i[22]
  PIN trng_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1496.000 631.490 1500.000 ;
    END
  END trng_wb_dat_i[23]
  PIN trng_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 1496.000 642.530 1500.000 ;
    END
  END trng_wb_dat_i[24]
  PIN trng_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 1496.000 646.670 1500.000 ;
    END
  END trng_wb_dat_i[25]
  PIN trng_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 685.480 1000.000 686.080 ;
    END
  END trng_wb_dat_i[26]
  PIN trng_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 738.520 1000.000 739.120 ;
    END
  END trng_wb_dat_i[27]
  PIN trng_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END trng_wb_dat_i[28]
  PIN trng_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 1496.000 665.070 1500.000 ;
    END
  END trng_wb_dat_i[29]
  PIN trng_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END trng_wb_dat_i[2]
  PIN trng_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 1496.000 676.110 1500.000 ;
    END
  END trng_wb_dat_i[30]
  PIN trng_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END trng_wb_dat_i[31]
  PIN trng_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 1496.000 464.970 1500.000 ;
    END
  END trng_wb_dat_i[3]
  PIN trng_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 142.840 1000.000 143.440 ;
    END
  END trng_wb_dat_i[4]
  PIN trng_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 1496.000 487.050 1500.000 ;
    END
  END trng_wb_dat_i[5]
  PIN trng_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END trng_wb_dat_i[6]
  PIN trng_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 1496.000 498.090 1500.000 ;
    END
  END trng_wb_dat_i[7]
  PIN trng_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 1496.000 509.590 1500.000 ;
    END
  END trng_wb_dat_i[8]
  PIN trng_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END trng_wb_dat_i[9]
  PIN trng_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 1496.000 442.890 1500.000 ;
    END
  END trng_wb_dat_o[0]
  PIN trng_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END trng_wb_dat_o[10]
  PIN trng_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END trng_wb_dat_o[11]
  PIN trng_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 387.640 1000.000 388.240 ;
    END
  END trng_wb_dat_o[12]
  PIN trng_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 408.720 1000.000 409.320 ;
    END
  END trng_wb_dat_o[13]
  PIN trng_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END trng_wb_dat_o[14]
  PIN trng_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 1496.000 557.430 1500.000 ;
    END
  END trng_wb_dat_o[15]
  PIN trng_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END trng_wb_dat_o[16]
  PIN trng_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 514.800 1000.000 515.400 ;
    END
  END trng_wb_dat_o[17]
  PIN trng_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END trng_wb_dat_o[18]
  PIN trng_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END trng_wb_dat_o[19]
  PIN trng_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END trng_wb_dat_o[1]
  PIN trng_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 546.760 1000.000 547.360 ;
    END
  END trng_wb_dat_o[20]
  PIN trng_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END trng_wb_dat_o[21]
  PIN trng_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END trng_wb_dat_o[22]
  PIN trng_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 1496.000 635.170 1500.000 ;
    END
  END trng_wb_dat_o[23]
  PIN trng_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 610.680 1000.000 611.280 ;
    END
  END trng_wb_dat_o[24]
  PIN trng_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END trng_wb_dat_o[25]
  PIN trng_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 1496.000 650.350 1500.000 ;
    END
  END trng_wb_dat_o[26]
  PIN trng_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END trng_wb_dat_o[27]
  PIN trng_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 770.480 1000.000 771.080 ;
    END
  END trng_wb_dat_o[28]
  PIN trng_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 823.520 1000.000 824.120 ;
    END
  END trng_wb_dat_o[29]
  PIN trng_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END trng_wb_dat_o[2]
  PIN trng_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 1496.000 679.790 1500.000 ;
    END
  END trng_wb_dat_o[30]
  PIN trng_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END trng_wb_dat_o[31]
  PIN trng_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 110.880 1000.000 111.480 ;
    END
  END trng_wb_dat_o[3]
  PIN trng_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END trng_wb_dat_o[4]
  PIN trng_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END trng_wb_dat_o[5]
  PIN trng_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 195.880 1000.000 196.480 ;
    END
  END trng_wb_dat_o[6]
  PIN trng_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 248.920 1000.000 249.520 ;
    END
  END trng_wb_dat_o[7]
  PIN trng_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END trng_wb_dat_o[8]
  PIN trng_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END trng_wb_dat_o[9]
  PIN trng_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END trng_wb_stb_o
  PIN trng_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 1496.000 427.710 1500.000 ;
    END
  END trng_wb_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 1487.925 ;
      LAYER met1 ;
        RECT 1.910 4.460 999.050 1488.080 ;
      LAYER met2 ;
        RECT 2.490 1495.720 5.330 1496.410 ;
        RECT 6.170 1495.720 9.010 1496.410 ;
        RECT 9.850 1495.720 12.690 1496.410 ;
        RECT 13.530 1495.720 16.370 1496.410 ;
        RECT 17.210 1495.720 20.050 1496.410 ;
        RECT 20.890 1495.720 23.730 1496.410 ;
        RECT 24.570 1495.720 27.410 1496.410 ;
        RECT 28.250 1495.720 31.090 1496.410 ;
        RECT 31.930 1495.720 34.770 1496.410 ;
        RECT 35.610 1495.720 38.450 1496.410 ;
        RECT 39.290 1495.720 42.130 1496.410 ;
        RECT 42.970 1495.720 45.810 1496.410 ;
        RECT 46.650 1495.720 49.490 1496.410 ;
        RECT 50.330 1495.720 53.170 1496.410 ;
        RECT 54.010 1495.720 56.850 1496.410 ;
        RECT 57.690 1495.720 60.530 1496.410 ;
        RECT 61.370 1495.720 64.210 1496.410 ;
        RECT 65.050 1495.720 67.890 1496.410 ;
        RECT 68.730 1495.720 71.570 1496.410 ;
        RECT 72.410 1495.720 75.710 1496.410 ;
        RECT 76.550 1495.720 79.390 1496.410 ;
        RECT 80.230 1495.720 83.070 1496.410 ;
        RECT 83.910 1495.720 86.750 1496.410 ;
        RECT 87.590 1495.720 90.430 1496.410 ;
        RECT 91.270 1495.720 94.110 1496.410 ;
        RECT 94.950 1495.720 97.790 1496.410 ;
        RECT 98.630 1495.720 101.470 1496.410 ;
        RECT 102.310 1495.720 105.150 1496.410 ;
        RECT 105.990 1495.720 108.830 1496.410 ;
        RECT 109.670 1495.720 112.510 1496.410 ;
        RECT 113.350 1495.720 116.190 1496.410 ;
        RECT 117.030 1495.720 119.870 1496.410 ;
        RECT 120.710 1495.720 123.550 1496.410 ;
        RECT 124.390 1495.720 127.230 1496.410 ;
        RECT 128.070 1495.720 130.910 1496.410 ;
        RECT 131.750 1495.720 134.590 1496.410 ;
        RECT 135.430 1495.720 138.270 1496.410 ;
        RECT 139.110 1495.720 141.950 1496.410 ;
        RECT 142.790 1495.720 146.090 1496.410 ;
        RECT 146.930 1495.720 149.770 1496.410 ;
        RECT 150.610 1495.720 153.450 1496.410 ;
        RECT 154.290 1495.720 157.130 1496.410 ;
        RECT 157.970 1495.720 160.810 1496.410 ;
        RECT 161.650 1495.720 164.490 1496.410 ;
        RECT 165.330 1495.720 168.170 1496.410 ;
        RECT 169.010 1495.720 171.850 1496.410 ;
        RECT 172.690 1495.720 175.530 1496.410 ;
        RECT 176.370 1495.720 179.210 1496.410 ;
        RECT 180.050 1495.720 182.890 1496.410 ;
        RECT 183.730 1495.720 186.570 1496.410 ;
        RECT 187.410 1495.720 190.250 1496.410 ;
        RECT 191.090 1495.720 193.930 1496.410 ;
        RECT 194.770 1495.720 197.610 1496.410 ;
        RECT 198.450 1495.720 201.290 1496.410 ;
        RECT 202.130 1495.720 204.970 1496.410 ;
        RECT 205.810 1495.720 208.650 1496.410 ;
        RECT 209.490 1495.720 212.330 1496.410 ;
        RECT 213.170 1495.720 216.470 1496.410 ;
        RECT 217.310 1495.720 220.150 1496.410 ;
        RECT 220.990 1495.720 223.830 1496.410 ;
        RECT 224.670 1495.720 227.510 1496.410 ;
        RECT 228.350 1495.720 231.190 1496.410 ;
        RECT 232.030 1495.720 234.870 1496.410 ;
        RECT 235.710 1495.720 238.550 1496.410 ;
        RECT 239.390 1495.720 242.230 1496.410 ;
        RECT 243.070 1495.720 245.910 1496.410 ;
        RECT 246.750 1495.720 249.590 1496.410 ;
        RECT 250.430 1495.720 253.270 1496.410 ;
        RECT 254.110 1495.720 256.950 1496.410 ;
        RECT 257.790 1495.720 260.630 1496.410 ;
        RECT 261.470 1495.720 264.310 1496.410 ;
        RECT 265.150 1495.720 267.990 1496.410 ;
        RECT 268.830 1495.720 271.670 1496.410 ;
        RECT 272.510 1495.720 275.350 1496.410 ;
        RECT 276.190 1495.720 279.030 1496.410 ;
        RECT 279.870 1495.720 282.710 1496.410 ;
        RECT 283.550 1495.720 286.390 1496.410 ;
        RECT 287.230 1495.720 290.530 1496.410 ;
        RECT 291.370 1495.720 294.210 1496.410 ;
        RECT 295.050 1495.720 297.890 1496.410 ;
        RECT 298.730 1495.720 301.570 1496.410 ;
        RECT 302.410 1495.720 305.250 1496.410 ;
        RECT 306.090 1495.720 308.930 1496.410 ;
        RECT 309.770 1495.720 312.610 1496.410 ;
        RECT 313.450 1495.720 316.290 1496.410 ;
        RECT 317.130 1495.720 319.970 1496.410 ;
        RECT 320.810 1495.720 323.650 1496.410 ;
        RECT 324.490 1495.720 327.330 1496.410 ;
        RECT 328.170 1495.720 331.010 1496.410 ;
        RECT 331.850 1495.720 334.690 1496.410 ;
        RECT 335.530 1495.720 338.370 1496.410 ;
        RECT 339.210 1495.720 342.050 1496.410 ;
        RECT 342.890 1495.720 345.730 1496.410 ;
        RECT 346.570 1495.720 349.410 1496.410 ;
        RECT 350.250 1495.720 353.090 1496.410 ;
        RECT 353.930 1495.720 356.770 1496.410 ;
        RECT 357.610 1495.720 360.910 1496.410 ;
        RECT 361.750 1495.720 364.590 1496.410 ;
        RECT 365.430 1495.720 368.270 1496.410 ;
        RECT 369.110 1495.720 371.950 1496.410 ;
        RECT 372.790 1495.720 375.630 1496.410 ;
        RECT 376.470 1495.720 379.310 1496.410 ;
        RECT 380.150 1495.720 382.990 1496.410 ;
        RECT 383.830 1495.720 386.670 1496.410 ;
        RECT 387.510 1495.720 390.350 1496.410 ;
        RECT 391.190 1495.720 394.030 1496.410 ;
        RECT 394.870 1495.720 397.710 1496.410 ;
        RECT 398.550 1495.720 401.390 1496.410 ;
        RECT 402.230 1495.720 405.070 1496.410 ;
        RECT 405.910 1495.720 408.750 1496.410 ;
        RECT 409.590 1495.720 412.430 1496.410 ;
        RECT 413.270 1495.720 416.110 1496.410 ;
        RECT 416.950 1495.720 419.790 1496.410 ;
        RECT 420.630 1495.720 423.470 1496.410 ;
        RECT 424.310 1495.720 427.150 1496.410 ;
        RECT 427.990 1495.720 431.290 1496.410 ;
        RECT 432.130 1495.720 434.970 1496.410 ;
        RECT 435.810 1495.720 438.650 1496.410 ;
        RECT 439.490 1495.720 442.330 1496.410 ;
        RECT 443.170 1495.720 446.010 1496.410 ;
        RECT 446.850 1495.720 449.690 1496.410 ;
        RECT 450.530 1495.720 453.370 1496.410 ;
        RECT 454.210 1495.720 457.050 1496.410 ;
        RECT 457.890 1495.720 460.730 1496.410 ;
        RECT 461.570 1495.720 464.410 1496.410 ;
        RECT 465.250 1495.720 468.090 1496.410 ;
        RECT 468.930 1495.720 471.770 1496.410 ;
        RECT 472.610 1495.720 475.450 1496.410 ;
        RECT 476.290 1495.720 479.130 1496.410 ;
        RECT 479.970 1495.720 482.810 1496.410 ;
        RECT 483.650 1495.720 486.490 1496.410 ;
        RECT 487.330 1495.720 490.170 1496.410 ;
        RECT 491.010 1495.720 493.850 1496.410 ;
        RECT 494.690 1495.720 497.530 1496.410 ;
        RECT 498.370 1495.720 501.670 1496.410 ;
        RECT 502.510 1495.720 505.350 1496.410 ;
        RECT 506.190 1495.720 509.030 1496.410 ;
        RECT 509.870 1495.720 512.710 1496.410 ;
        RECT 513.550 1495.720 516.390 1496.410 ;
        RECT 517.230 1495.720 520.070 1496.410 ;
        RECT 520.910 1495.720 523.750 1496.410 ;
        RECT 524.590 1495.720 527.430 1496.410 ;
        RECT 528.270 1495.720 531.110 1496.410 ;
        RECT 531.950 1495.720 534.790 1496.410 ;
        RECT 535.630 1495.720 538.470 1496.410 ;
        RECT 539.310 1495.720 542.150 1496.410 ;
        RECT 542.990 1495.720 545.830 1496.410 ;
        RECT 546.670 1495.720 549.510 1496.410 ;
        RECT 550.350 1495.720 553.190 1496.410 ;
        RECT 554.030 1495.720 556.870 1496.410 ;
        RECT 557.710 1495.720 560.550 1496.410 ;
        RECT 561.390 1495.720 564.230 1496.410 ;
        RECT 565.070 1495.720 567.910 1496.410 ;
        RECT 568.750 1495.720 571.590 1496.410 ;
        RECT 572.430 1495.720 575.730 1496.410 ;
        RECT 576.570 1495.720 579.410 1496.410 ;
        RECT 580.250 1495.720 583.090 1496.410 ;
        RECT 583.930 1495.720 586.770 1496.410 ;
        RECT 587.610 1495.720 590.450 1496.410 ;
        RECT 591.290 1495.720 594.130 1496.410 ;
        RECT 594.970 1495.720 597.810 1496.410 ;
        RECT 598.650 1495.720 601.490 1496.410 ;
        RECT 602.330 1495.720 605.170 1496.410 ;
        RECT 606.010 1495.720 608.850 1496.410 ;
        RECT 609.690 1495.720 612.530 1496.410 ;
        RECT 613.370 1495.720 616.210 1496.410 ;
        RECT 617.050 1495.720 619.890 1496.410 ;
        RECT 620.730 1495.720 623.570 1496.410 ;
        RECT 624.410 1495.720 627.250 1496.410 ;
        RECT 628.090 1495.720 630.930 1496.410 ;
        RECT 631.770 1495.720 634.610 1496.410 ;
        RECT 635.450 1495.720 638.290 1496.410 ;
        RECT 639.130 1495.720 641.970 1496.410 ;
        RECT 642.810 1495.720 646.110 1496.410 ;
        RECT 646.950 1495.720 649.790 1496.410 ;
        RECT 650.630 1495.720 653.470 1496.410 ;
        RECT 654.310 1495.720 657.150 1496.410 ;
        RECT 657.990 1495.720 660.830 1496.410 ;
        RECT 661.670 1495.720 664.510 1496.410 ;
        RECT 665.350 1495.720 668.190 1496.410 ;
        RECT 669.030 1495.720 671.870 1496.410 ;
        RECT 672.710 1495.720 675.550 1496.410 ;
        RECT 676.390 1495.720 679.230 1496.410 ;
        RECT 680.070 1495.720 682.910 1496.410 ;
        RECT 683.750 1495.720 686.590 1496.410 ;
        RECT 687.430 1495.720 690.270 1496.410 ;
        RECT 691.110 1495.720 693.950 1496.410 ;
        RECT 694.790 1495.720 697.630 1496.410 ;
        RECT 698.470 1495.720 701.310 1496.410 ;
        RECT 702.150 1495.720 704.990 1496.410 ;
        RECT 705.830 1495.720 708.670 1496.410 ;
        RECT 709.510 1495.720 712.350 1496.410 ;
        RECT 713.190 1495.720 716.490 1496.410 ;
        RECT 717.330 1495.720 720.170 1496.410 ;
        RECT 721.010 1495.720 723.850 1496.410 ;
        RECT 724.690 1495.720 727.530 1496.410 ;
        RECT 728.370 1495.720 731.210 1496.410 ;
        RECT 732.050 1495.720 734.890 1496.410 ;
        RECT 735.730 1495.720 738.570 1496.410 ;
        RECT 739.410 1495.720 742.250 1496.410 ;
        RECT 743.090 1495.720 745.930 1496.410 ;
        RECT 746.770 1495.720 749.610 1496.410 ;
        RECT 750.450 1495.720 753.290 1496.410 ;
        RECT 754.130 1495.720 756.970 1496.410 ;
        RECT 757.810 1495.720 760.650 1496.410 ;
        RECT 761.490 1495.720 764.330 1496.410 ;
        RECT 765.170 1495.720 768.010 1496.410 ;
        RECT 768.850 1495.720 771.690 1496.410 ;
        RECT 772.530 1495.720 775.370 1496.410 ;
        RECT 776.210 1495.720 779.050 1496.410 ;
        RECT 779.890 1495.720 782.730 1496.410 ;
        RECT 783.570 1495.720 786.410 1496.410 ;
        RECT 787.250 1495.720 790.550 1496.410 ;
        RECT 791.390 1495.720 794.230 1496.410 ;
        RECT 795.070 1495.720 797.910 1496.410 ;
        RECT 798.750 1495.720 801.590 1496.410 ;
        RECT 802.430 1495.720 805.270 1496.410 ;
        RECT 806.110 1495.720 808.950 1496.410 ;
        RECT 809.790 1495.720 812.630 1496.410 ;
        RECT 813.470 1495.720 816.310 1496.410 ;
        RECT 817.150 1495.720 819.990 1496.410 ;
        RECT 820.830 1495.720 823.670 1496.410 ;
        RECT 824.510 1495.720 827.350 1496.410 ;
        RECT 828.190 1495.720 831.030 1496.410 ;
        RECT 831.870 1495.720 834.710 1496.410 ;
        RECT 835.550 1495.720 838.390 1496.410 ;
        RECT 839.230 1495.720 842.070 1496.410 ;
        RECT 842.910 1495.720 845.750 1496.410 ;
        RECT 846.590 1495.720 849.430 1496.410 ;
        RECT 850.270 1495.720 853.110 1496.410 ;
        RECT 853.950 1495.720 856.790 1496.410 ;
        RECT 857.630 1495.720 860.930 1496.410 ;
        RECT 861.770 1495.720 864.610 1496.410 ;
        RECT 865.450 1495.720 868.290 1496.410 ;
        RECT 869.130 1495.720 871.970 1496.410 ;
        RECT 872.810 1495.720 875.650 1496.410 ;
        RECT 876.490 1495.720 879.330 1496.410 ;
        RECT 880.170 1495.720 883.010 1496.410 ;
        RECT 883.850 1495.720 886.690 1496.410 ;
        RECT 887.530 1495.720 890.370 1496.410 ;
        RECT 891.210 1495.720 894.050 1496.410 ;
        RECT 894.890 1495.720 897.730 1496.410 ;
        RECT 898.570 1495.720 901.410 1496.410 ;
        RECT 902.250 1495.720 905.090 1496.410 ;
        RECT 905.930 1495.720 908.770 1496.410 ;
        RECT 909.610 1495.720 912.450 1496.410 ;
        RECT 913.290 1495.720 916.130 1496.410 ;
        RECT 916.970 1495.720 919.810 1496.410 ;
        RECT 920.650 1495.720 923.490 1496.410 ;
        RECT 924.330 1495.720 927.170 1496.410 ;
        RECT 928.010 1495.720 931.310 1496.410 ;
        RECT 932.150 1495.720 934.990 1496.410 ;
        RECT 935.830 1495.720 938.670 1496.410 ;
        RECT 939.510 1495.720 942.350 1496.410 ;
        RECT 943.190 1495.720 946.030 1496.410 ;
        RECT 946.870 1495.720 949.710 1496.410 ;
        RECT 950.550 1495.720 953.390 1496.410 ;
        RECT 954.230 1495.720 957.070 1496.410 ;
        RECT 957.910 1495.720 960.750 1496.410 ;
        RECT 961.590 1495.720 964.430 1496.410 ;
        RECT 965.270 1495.720 968.110 1496.410 ;
        RECT 968.950 1495.720 971.790 1496.410 ;
        RECT 972.630 1495.720 975.470 1496.410 ;
        RECT 976.310 1495.720 979.150 1496.410 ;
        RECT 979.990 1495.720 982.830 1496.410 ;
        RECT 983.670 1495.720 986.510 1496.410 ;
        RECT 987.350 1495.720 990.190 1496.410 ;
        RECT 991.030 1495.720 993.870 1496.410 ;
        RECT 994.710 1495.720 997.550 1496.410 ;
        RECT 998.390 1495.720 999.020 1496.410 ;
        RECT 1.940 4.280 999.020 1495.720 ;
        RECT 2.490 3.670 5.330 4.280 ;
        RECT 6.170 3.670 9.470 4.280 ;
        RECT 10.310 3.670 13.610 4.280 ;
        RECT 14.450 3.670 17.750 4.280 ;
        RECT 18.590 3.670 21.890 4.280 ;
        RECT 22.730 3.670 26.030 4.280 ;
        RECT 26.870 3.670 30.170 4.280 ;
        RECT 31.010 3.670 33.850 4.280 ;
        RECT 34.690 3.670 37.990 4.280 ;
        RECT 38.830 3.670 42.130 4.280 ;
        RECT 42.970 3.670 46.270 4.280 ;
        RECT 47.110 3.670 50.410 4.280 ;
        RECT 51.250 3.670 54.550 4.280 ;
        RECT 55.390 3.670 58.690 4.280 ;
        RECT 59.530 3.670 62.830 4.280 ;
        RECT 63.670 3.670 66.510 4.280 ;
        RECT 67.350 3.670 70.650 4.280 ;
        RECT 71.490 3.670 74.790 4.280 ;
        RECT 75.630 3.670 78.930 4.280 ;
        RECT 79.770 3.670 83.070 4.280 ;
        RECT 83.910 3.670 87.210 4.280 ;
        RECT 88.050 3.670 91.350 4.280 ;
        RECT 92.190 3.670 95.490 4.280 ;
        RECT 96.330 3.670 99.170 4.280 ;
        RECT 100.010 3.670 103.310 4.280 ;
        RECT 104.150 3.670 107.450 4.280 ;
        RECT 108.290 3.670 111.590 4.280 ;
        RECT 112.430 3.670 115.730 4.280 ;
        RECT 116.570 3.670 119.870 4.280 ;
        RECT 120.710 3.670 124.010 4.280 ;
        RECT 124.850 3.670 128.150 4.280 ;
        RECT 128.990 3.670 131.830 4.280 ;
        RECT 132.670 3.670 135.970 4.280 ;
        RECT 136.810 3.670 140.110 4.280 ;
        RECT 140.950 3.670 144.250 4.280 ;
        RECT 145.090 3.670 148.390 4.280 ;
        RECT 149.230 3.670 152.530 4.280 ;
        RECT 153.370 3.670 156.670 4.280 ;
        RECT 157.510 3.670 160.810 4.280 ;
        RECT 161.650 3.670 164.490 4.280 ;
        RECT 165.330 3.670 168.630 4.280 ;
        RECT 169.470 3.670 172.770 4.280 ;
        RECT 173.610 3.670 176.910 4.280 ;
        RECT 177.750 3.670 181.050 4.280 ;
        RECT 181.890 3.670 185.190 4.280 ;
        RECT 186.030 3.670 189.330 4.280 ;
        RECT 190.170 3.670 193.470 4.280 ;
        RECT 194.310 3.670 197.150 4.280 ;
        RECT 197.990 3.670 201.290 4.280 ;
        RECT 202.130 3.670 205.430 4.280 ;
        RECT 206.270 3.670 209.570 4.280 ;
        RECT 210.410 3.670 213.710 4.280 ;
        RECT 214.550 3.670 217.850 4.280 ;
        RECT 218.690 3.670 221.990 4.280 ;
        RECT 222.830 3.670 226.130 4.280 ;
        RECT 226.970 3.670 229.810 4.280 ;
        RECT 230.650 3.670 233.950 4.280 ;
        RECT 234.790 3.670 238.090 4.280 ;
        RECT 238.930 3.670 242.230 4.280 ;
        RECT 243.070 3.670 246.370 4.280 ;
        RECT 247.210 3.670 250.510 4.280 ;
        RECT 251.350 3.670 254.650 4.280 ;
        RECT 255.490 3.670 258.790 4.280 ;
        RECT 259.630 3.670 262.470 4.280 ;
        RECT 263.310 3.670 266.610 4.280 ;
        RECT 267.450 3.670 270.750 4.280 ;
        RECT 271.590 3.670 274.890 4.280 ;
        RECT 275.730 3.670 279.030 4.280 ;
        RECT 279.870 3.670 283.170 4.280 ;
        RECT 284.010 3.670 287.310 4.280 ;
        RECT 288.150 3.670 291.450 4.280 ;
        RECT 292.290 3.670 295.130 4.280 ;
        RECT 295.970 3.670 299.270 4.280 ;
        RECT 300.110 3.670 303.410 4.280 ;
        RECT 304.250 3.670 307.550 4.280 ;
        RECT 308.390 3.670 311.690 4.280 ;
        RECT 312.530 3.670 315.830 4.280 ;
        RECT 316.670 3.670 319.970 4.280 ;
        RECT 320.810 3.670 324.110 4.280 ;
        RECT 324.950 3.670 327.790 4.280 ;
        RECT 328.630 3.670 331.930 4.280 ;
        RECT 332.770 3.670 336.070 4.280 ;
        RECT 336.910 3.670 340.210 4.280 ;
        RECT 341.050 3.670 344.350 4.280 ;
        RECT 345.190 3.670 348.490 4.280 ;
        RECT 349.330 3.670 352.630 4.280 ;
        RECT 353.470 3.670 356.310 4.280 ;
        RECT 357.150 3.670 360.450 4.280 ;
        RECT 361.290 3.670 364.590 4.280 ;
        RECT 365.430 3.670 368.730 4.280 ;
        RECT 369.570 3.670 372.870 4.280 ;
        RECT 373.710 3.670 377.010 4.280 ;
        RECT 377.850 3.670 381.150 4.280 ;
        RECT 381.990 3.670 385.290 4.280 ;
        RECT 386.130 3.670 388.970 4.280 ;
        RECT 389.810 3.670 393.110 4.280 ;
        RECT 393.950 3.670 397.250 4.280 ;
        RECT 398.090 3.670 401.390 4.280 ;
        RECT 402.230 3.670 405.530 4.280 ;
        RECT 406.370 3.670 409.670 4.280 ;
        RECT 410.510 3.670 413.810 4.280 ;
        RECT 414.650 3.670 417.950 4.280 ;
        RECT 418.790 3.670 421.630 4.280 ;
        RECT 422.470 3.670 425.770 4.280 ;
        RECT 426.610 3.670 429.910 4.280 ;
        RECT 430.750 3.670 434.050 4.280 ;
        RECT 434.890 3.670 438.190 4.280 ;
        RECT 439.030 3.670 442.330 4.280 ;
        RECT 443.170 3.670 446.470 4.280 ;
        RECT 447.310 3.670 450.610 4.280 ;
        RECT 451.450 3.670 454.290 4.280 ;
        RECT 455.130 3.670 458.430 4.280 ;
        RECT 459.270 3.670 462.570 4.280 ;
        RECT 463.410 3.670 466.710 4.280 ;
        RECT 467.550 3.670 470.850 4.280 ;
        RECT 471.690 3.670 474.990 4.280 ;
        RECT 475.830 3.670 479.130 4.280 ;
        RECT 479.970 3.670 483.270 4.280 ;
        RECT 484.110 3.670 486.950 4.280 ;
        RECT 487.790 3.670 491.090 4.280 ;
        RECT 491.930 3.670 495.230 4.280 ;
        RECT 496.070 3.670 499.370 4.280 ;
        RECT 500.210 3.670 503.510 4.280 ;
        RECT 504.350 3.670 507.650 4.280 ;
        RECT 508.490 3.670 511.790 4.280 ;
        RECT 512.630 3.670 515.930 4.280 ;
        RECT 516.770 3.670 519.610 4.280 ;
        RECT 520.450 3.670 523.750 4.280 ;
        RECT 524.590 3.670 527.890 4.280 ;
        RECT 528.730 3.670 532.030 4.280 ;
        RECT 532.870 3.670 536.170 4.280 ;
        RECT 537.010 3.670 540.310 4.280 ;
        RECT 541.150 3.670 544.450 4.280 ;
        RECT 545.290 3.670 548.590 4.280 ;
        RECT 549.430 3.670 552.270 4.280 ;
        RECT 553.110 3.670 556.410 4.280 ;
        RECT 557.250 3.670 560.550 4.280 ;
        RECT 561.390 3.670 564.690 4.280 ;
        RECT 565.530 3.670 568.830 4.280 ;
        RECT 569.670 3.670 572.970 4.280 ;
        RECT 573.810 3.670 577.110 4.280 ;
        RECT 577.950 3.670 581.250 4.280 ;
        RECT 582.090 3.670 584.930 4.280 ;
        RECT 585.770 3.670 589.070 4.280 ;
        RECT 589.910 3.670 593.210 4.280 ;
        RECT 594.050 3.670 597.350 4.280 ;
        RECT 598.190 3.670 601.490 4.280 ;
        RECT 602.330 3.670 605.630 4.280 ;
        RECT 606.470 3.670 609.770 4.280 ;
        RECT 610.610 3.670 613.910 4.280 ;
        RECT 614.750 3.670 617.590 4.280 ;
        RECT 618.430 3.670 621.730 4.280 ;
        RECT 622.570 3.670 625.870 4.280 ;
        RECT 626.710 3.670 630.010 4.280 ;
        RECT 630.850 3.670 634.150 4.280 ;
        RECT 634.990 3.670 638.290 4.280 ;
        RECT 639.130 3.670 642.430 4.280 ;
        RECT 643.270 3.670 646.570 4.280 ;
        RECT 647.410 3.670 650.250 4.280 ;
        RECT 651.090 3.670 654.390 4.280 ;
        RECT 655.230 3.670 658.530 4.280 ;
        RECT 659.370 3.670 662.670 4.280 ;
        RECT 663.510 3.670 666.810 4.280 ;
        RECT 667.650 3.670 670.950 4.280 ;
        RECT 671.790 3.670 675.090 4.280 ;
        RECT 675.930 3.670 678.770 4.280 ;
        RECT 679.610 3.670 682.910 4.280 ;
        RECT 683.750 3.670 687.050 4.280 ;
        RECT 687.890 3.670 691.190 4.280 ;
        RECT 692.030 3.670 695.330 4.280 ;
        RECT 696.170 3.670 699.470 4.280 ;
        RECT 700.310 3.670 703.610 4.280 ;
        RECT 704.450 3.670 707.750 4.280 ;
        RECT 708.590 3.670 711.430 4.280 ;
        RECT 712.270 3.670 715.570 4.280 ;
        RECT 716.410 3.670 719.710 4.280 ;
        RECT 720.550 3.670 723.850 4.280 ;
        RECT 724.690 3.670 727.990 4.280 ;
        RECT 728.830 3.670 732.130 4.280 ;
        RECT 732.970 3.670 736.270 4.280 ;
        RECT 737.110 3.670 740.410 4.280 ;
        RECT 741.250 3.670 744.090 4.280 ;
        RECT 744.930 3.670 748.230 4.280 ;
        RECT 749.070 3.670 752.370 4.280 ;
        RECT 753.210 3.670 756.510 4.280 ;
        RECT 757.350 3.670 760.650 4.280 ;
        RECT 761.490 3.670 764.790 4.280 ;
        RECT 765.630 3.670 768.930 4.280 ;
        RECT 769.770 3.670 773.070 4.280 ;
        RECT 773.910 3.670 776.750 4.280 ;
        RECT 777.590 3.670 780.890 4.280 ;
        RECT 781.730 3.670 785.030 4.280 ;
        RECT 785.870 3.670 789.170 4.280 ;
        RECT 790.010 3.670 793.310 4.280 ;
        RECT 794.150 3.670 797.450 4.280 ;
        RECT 798.290 3.670 801.590 4.280 ;
        RECT 802.430 3.670 805.730 4.280 ;
        RECT 806.570 3.670 809.410 4.280 ;
        RECT 810.250 3.670 813.550 4.280 ;
        RECT 814.390 3.670 817.690 4.280 ;
        RECT 818.530 3.670 821.830 4.280 ;
        RECT 822.670 3.670 825.970 4.280 ;
        RECT 826.810 3.670 830.110 4.280 ;
        RECT 830.950 3.670 834.250 4.280 ;
        RECT 835.090 3.670 838.390 4.280 ;
        RECT 839.230 3.670 842.070 4.280 ;
        RECT 842.910 3.670 846.210 4.280 ;
        RECT 847.050 3.670 850.350 4.280 ;
        RECT 851.190 3.670 854.490 4.280 ;
        RECT 855.330 3.670 858.630 4.280 ;
        RECT 859.470 3.670 862.770 4.280 ;
        RECT 863.610 3.670 866.910 4.280 ;
        RECT 867.750 3.670 871.050 4.280 ;
        RECT 871.890 3.670 874.730 4.280 ;
        RECT 875.570 3.670 878.870 4.280 ;
        RECT 879.710 3.670 883.010 4.280 ;
        RECT 883.850 3.670 887.150 4.280 ;
        RECT 887.990 3.670 891.290 4.280 ;
        RECT 892.130 3.670 895.430 4.280 ;
        RECT 896.270 3.670 899.570 4.280 ;
        RECT 900.410 3.670 903.710 4.280 ;
        RECT 904.550 3.670 907.390 4.280 ;
        RECT 908.230 3.670 911.530 4.280 ;
        RECT 912.370 3.670 915.670 4.280 ;
        RECT 916.510 3.670 919.810 4.280 ;
        RECT 920.650 3.670 923.950 4.280 ;
        RECT 924.790 3.670 928.090 4.280 ;
        RECT 928.930 3.670 932.230 4.280 ;
        RECT 933.070 3.670 936.370 4.280 ;
        RECT 937.210 3.670 940.050 4.280 ;
        RECT 940.890 3.670 944.190 4.280 ;
        RECT 945.030 3.670 948.330 4.280 ;
        RECT 949.170 3.670 952.470 4.280 ;
        RECT 953.310 3.670 956.610 4.280 ;
        RECT 957.450 3.670 960.750 4.280 ;
        RECT 961.590 3.670 964.890 4.280 ;
        RECT 965.730 3.670 969.030 4.280 ;
        RECT 969.870 3.670 972.710 4.280 ;
        RECT 973.550 3.670 976.850 4.280 ;
        RECT 977.690 3.670 980.990 4.280 ;
        RECT 981.830 3.670 985.130 4.280 ;
        RECT 985.970 3.670 989.270 4.280 ;
        RECT 990.110 3.670 993.410 4.280 ;
        RECT 994.250 3.670 997.550 4.280 ;
        RECT 998.390 3.670 999.020 4.280 ;
      LAYER met3 ;
        RECT 4.400 1495.000 996.000 1495.145 ;
        RECT 4.400 1494.280 995.600 1495.000 ;
        RECT 4.000 1493.600 995.600 1494.280 ;
        RECT 4.000 1485.480 996.000 1493.600 ;
        RECT 4.400 1484.120 996.000 1485.480 ;
        RECT 4.400 1484.080 995.600 1484.120 ;
        RECT 4.000 1482.720 995.600 1484.080 ;
        RECT 4.000 1475.280 996.000 1482.720 ;
        RECT 4.400 1473.920 996.000 1475.280 ;
        RECT 4.400 1473.880 995.600 1473.920 ;
        RECT 4.000 1472.520 995.600 1473.880 ;
        RECT 4.000 1465.080 996.000 1472.520 ;
        RECT 4.400 1463.680 996.000 1465.080 ;
        RECT 4.000 1463.040 996.000 1463.680 ;
        RECT 4.000 1461.640 995.600 1463.040 ;
        RECT 4.000 1454.880 996.000 1461.640 ;
        RECT 4.400 1453.480 996.000 1454.880 ;
        RECT 4.000 1452.160 996.000 1453.480 ;
        RECT 4.000 1450.760 995.600 1452.160 ;
        RECT 4.000 1445.360 996.000 1450.760 ;
        RECT 4.400 1443.960 996.000 1445.360 ;
        RECT 4.000 1441.960 996.000 1443.960 ;
        RECT 4.000 1440.560 995.600 1441.960 ;
        RECT 4.000 1435.160 996.000 1440.560 ;
        RECT 4.400 1433.760 996.000 1435.160 ;
        RECT 4.000 1431.080 996.000 1433.760 ;
        RECT 4.000 1429.680 995.600 1431.080 ;
        RECT 4.000 1424.960 996.000 1429.680 ;
        RECT 4.400 1423.560 996.000 1424.960 ;
        RECT 4.000 1420.200 996.000 1423.560 ;
        RECT 4.000 1418.800 995.600 1420.200 ;
        RECT 4.000 1414.760 996.000 1418.800 ;
        RECT 4.400 1413.360 996.000 1414.760 ;
        RECT 4.000 1410.000 996.000 1413.360 ;
        RECT 4.000 1408.600 995.600 1410.000 ;
        RECT 4.000 1404.560 996.000 1408.600 ;
        RECT 4.400 1403.160 996.000 1404.560 ;
        RECT 4.000 1399.120 996.000 1403.160 ;
        RECT 4.000 1397.720 995.600 1399.120 ;
        RECT 4.000 1395.040 996.000 1397.720 ;
        RECT 4.400 1393.640 996.000 1395.040 ;
        RECT 4.000 1388.240 996.000 1393.640 ;
        RECT 4.000 1386.840 995.600 1388.240 ;
        RECT 4.000 1384.840 996.000 1386.840 ;
        RECT 4.400 1383.440 996.000 1384.840 ;
        RECT 4.000 1378.040 996.000 1383.440 ;
        RECT 4.000 1376.640 995.600 1378.040 ;
        RECT 4.000 1374.640 996.000 1376.640 ;
        RECT 4.400 1373.240 996.000 1374.640 ;
        RECT 4.000 1367.160 996.000 1373.240 ;
        RECT 4.000 1365.760 995.600 1367.160 ;
        RECT 4.000 1364.440 996.000 1365.760 ;
        RECT 4.400 1363.040 996.000 1364.440 ;
        RECT 4.000 1356.280 996.000 1363.040 ;
        RECT 4.000 1354.880 995.600 1356.280 ;
        RECT 4.000 1354.240 996.000 1354.880 ;
        RECT 4.400 1352.840 996.000 1354.240 ;
        RECT 4.000 1346.080 996.000 1352.840 ;
        RECT 4.000 1344.720 995.600 1346.080 ;
        RECT 4.400 1344.680 995.600 1344.720 ;
        RECT 4.400 1343.320 996.000 1344.680 ;
        RECT 4.000 1335.200 996.000 1343.320 ;
        RECT 4.000 1334.520 995.600 1335.200 ;
        RECT 4.400 1333.800 995.600 1334.520 ;
        RECT 4.400 1333.120 996.000 1333.800 ;
        RECT 4.000 1325.000 996.000 1333.120 ;
        RECT 4.000 1324.320 995.600 1325.000 ;
        RECT 4.400 1323.600 995.600 1324.320 ;
        RECT 4.400 1322.920 996.000 1323.600 ;
        RECT 4.000 1314.120 996.000 1322.920 ;
        RECT 4.400 1312.720 995.600 1314.120 ;
        RECT 4.000 1303.920 996.000 1312.720 ;
        RECT 4.400 1303.240 996.000 1303.920 ;
        RECT 4.400 1302.520 995.600 1303.240 ;
        RECT 4.000 1301.840 995.600 1302.520 ;
        RECT 4.000 1294.400 996.000 1301.840 ;
        RECT 4.400 1293.040 996.000 1294.400 ;
        RECT 4.400 1293.000 995.600 1293.040 ;
        RECT 4.000 1291.640 995.600 1293.000 ;
        RECT 4.000 1284.200 996.000 1291.640 ;
        RECT 4.400 1282.800 996.000 1284.200 ;
        RECT 4.000 1282.160 996.000 1282.800 ;
        RECT 4.000 1280.760 995.600 1282.160 ;
        RECT 4.000 1274.000 996.000 1280.760 ;
        RECT 4.400 1272.600 996.000 1274.000 ;
        RECT 4.000 1271.280 996.000 1272.600 ;
        RECT 4.000 1269.880 995.600 1271.280 ;
        RECT 4.000 1263.800 996.000 1269.880 ;
        RECT 4.400 1262.400 996.000 1263.800 ;
        RECT 4.000 1261.080 996.000 1262.400 ;
        RECT 4.000 1259.680 995.600 1261.080 ;
        RECT 4.000 1253.600 996.000 1259.680 ;
        RECT 4.400 1252.200 996.000 1253.600 ;
        RECT 4.000 1250.200 996.000 1252.200 ;
        RECT 4.000 1248.800 995.600 1250.200 ;
        RECT 4.000 1244.080 996.000 1248.800 ;
        RECT 4.400 1242.680 996.000 1244.080 ;
        RECT 4.000 1239.320 996.000 1242.680 ;
        RECT 4.000 1237.920 995.600 1239.320 ;
        RECT 4.000 1233.880 996.000 1237.920 ;
        RECT 4.400 1232.480 996.000 1233.880 ;
        RECT 4.000 1229.120 996.000 1232.480 ;
        RECT 4.000 1227.720 995.600 1229.120 ;
        RECT 4.000 1223.680 996.000 1227.720 ;
        RECT 4.400 1222.280 996.000 1223.680 ;
        RECT 4.000 1218.240 996.000 1222.280 ;
        RECT 4.000 1216.840 995.600 1218.240 ;
        RECT 4.000 1213.480 996.000 1216.840 ;
        RECT 4.400 1212.080 996.000 1213.480 ;
        RECT 4.000 1207.360 996.000 1212.080 ;
        RECT 4.000 1205.960 995.600 1207.360 ;
        RECT 4.000 1203.280 996.000 1205.960 ;
        RECT 4.400 1201.880 996.000 1203.280 ;
        RECT 4.000 1197.160 996.000 1201.880 ;
        RECT 4.000 1195.760 995.600 1197.160 ;
        RECT 4.000 1193.760 996.000 1195.760 ;
        RECT 4.400 1192.360 996.000 1193.760 ;
        RECT 4.000 1186.280 996.000 1192.360 ;
        RECT 4.000 1184.880 995.600 1186.280 ;
        RECT 4.000 1183.560 996.000 1184.880 ;
        RECT 4.400 1182.160 996.000 1183.560 ;
        RECT 4.000 1175.400 996.000 1182.160 ;
        RECT 4.000 1174.000 995.600 1175.400 ;
        RECT 4.000 1173.360 996.000 1174.000 ;
        RECT 4.400 1171.960 996.000 1173.360 ;
        RECT 4.000 1165.200 996.000 1171.960 ;
        RECT 4.000 1163.800 995.600 1165.200 ;
        RECT 4.000 1163.160 996.000 1163.800 ;
        RECT 4.400 1161.760 996.000 1163.160 ;
        RECT 4.000 1154.320 996.000 1161.760 ;
        RECT 4.000 1152.960 995.600 1154.320 ;
        RECT 4.400 1152.920 995.600 1152.960 ;
        RECT 4.400 1151.560 996.000 1152.920 ;
        RECT 4.000 1144.120 996.000 1151.560 ;
        RECT 4.000 1143.440 995.600 1144.120 ;
        RECT 4.400 1142.720 995.600 1143.440 ;
        RECT 4.400 1142.040 996.000 1142.720 ;
        RECT 4.000 1133.240 996.000 1142.040 ;
        RECT 4.400 1131.840 995.600 1133.240 ;
        RECT 4.000 1123.040 996.000 1131.840 ;
        RECT 4.400 1122.360 996.000 1123.040 ;
        RECT 4.400 1121.640 995.600 1122.360 ;
        RECT 4.000 1120.960 995.600 1121.640 ;
        RECT 4.000 1112.840 996.000 1120.960 ;
        RECT 4.400 1112.160 996.000 1112.840 ;
        RECT 4.400 1111.440 995.600 1112.160 ;
        RECT 4.000 1110.760 995.600 1111.440 ;
        RECT 4.000 1102.640 996.000 1110.760 ;
        RECT 4.400 1101.280 996.000 1102.640 ;
        RECT 4.400 1101.240 995.600 1101.280 ;
        RECT 4.000 1099.880 995.600 1101.240 ;
        RECT 4.000 1092.440 996.000 1099.880 ;
        RECT 4.400 1091.040 996.000 1092.440 ;
        RECT 4.000 1090.400 996.000 1091.040 ;
        RECT 4.000 1089.000 995.600 1090.400 ;
        RECT 4.000 1082.920 996.000 1089.000 ;
        RECT 4.400 1081.520 996.000 1082.920 ;
        RECT 4.000 1080.200 996.000 1081.520 ;
        RECT 4.000 1078.800 995.600 1080.200 ;
        RECT 4.000 1072.720 996.000 1078.800 ;
        RECT 4.400 1071.320 996.000 1072.720 ;
        RECT 4.000 1069.320 996.000 1071.320 ;
        RECT 4.000 1067.920 995.600 1069.320 ;
        RECT 4.000 1062.520 996.000 1067.920 ;
        RECT 4.400 1061.120 996.000 1062.520 ;
        RECT 4.000 1058.440 996.000 1061.120 ;
        RECT 4.000 1057.040 995.600 1058.440 ;
        RECT 4.000 1052.320 996.000 1057.040 ;
        RECT 4.400 1050.920 996.000 1052.320 ;
        RECT 4.000 1048.240 996.000 1050.920 ;
        RECT 4.000 1046.840 995.600 1048.240 ;
        RECT 4.000 1042.120 996.000 1046.840 ;
        RECT 4.400 1040.720 996.000 1042.120 ;
        RECT 4.000 1037.360 996.000 1040.720 ;
        RECT 4.000 1035.960 995.600 1037.360 ;
        RECT 4.000 1032.600 996.000 1035.960 ;
        RECT 4.400 1031.200 996.000 1032.600 ;
        RECT 4.000 1026.480 996.000 1031.200 ;
        RECT 4.000 1025.080 995.600 1026.480 ;
        RECT 4.000 1022.400 996.000 1025.080 ;
        RECT 4.400 1021.000 996.000 1022.400 ;
        RECT 4.000 1016.280 996.000 1021.000 ;
        RECT 4.000 1014.880 995.600 1016.280 ;
        RECT 4.000 1012.200 996.000 1014.880 ;
        RECT 4.400 1010.800 996.000 1012.200 ;
        RECT 4.000 1005.400 996.000 1010.800 ;
        RECT 4.000 1004.000 995.600 1005.400 ;
        RECT 4.000 1002.000 996.000 1004.000 ;
        RECT 4.400 1000.600 996.000 1002.000 ;
        RECT 4.000 995.200 996.000 1000.600 ;
        RECT 4.000 993.800 995.600 995.200 ;
        RECT 4.000 991.800 996.000 993.800 ;
        RECT 4.400 990.400 996.000 991.800 ;
        RECT 4.000 984.320 996.000 990.400 ;
        RECT 4.000 982.920 995.600 984.320 ;
        RECT 4.000 982.280 996.000 982.920 ;
        RECT 4.400 980.880 996.000 982.280 ;
        RECT 4.000 973.440 996.000 980.880 ;
        RECT 4.000 972.080 995.600 973.440 ;
        RECT 4.400 972.040 995.600 972.080 ;
        RECT 4.400 970.680 996.000 972.040 ;
        RECT 4.000 963.240 996.000 970.680 ;
        RECT 4.000 961.880 995.600 963.240 ;
        RECT 4.400 961.840 995.600 961.880 ;
        RECT 4.400 960.480 996.000 961.840 ;
        RECT 4.000 952.360 996.000 960.480 ;
        RECT 4.000 951.680 995.600 952.360 ;
        RECT 4.400 950.960 995.600 951.680 ;
        RECT 4.400 950.280 996.000 950.960 ;
        RECT 4.000 941.480 996.000 950.280 ;
        RECT 4.400 940.080 995.600 941.480 ;
        RECT 4.000 931.960 996.000 940.080 ;
        RECT 4.400 931.280 996.000 931.960 ;
        RECT 4.400 930.560 995.600 931.280 ;
        RECT 4.000 929.880 995.600 930.560 ;
        RECT 4.000 921.760 996.000 929.880 ;
        RECT 4.400 920.400 996.000 921.760 ;
        RECT 4.400 920.360 995.600 920.400 ;
        RECT 4.000 919.000 995.600 920.360 ;
        RECT 4.000 911.560 996.000 919.000 ;
        RECT 4.400 910.160 996.000 911.560 ;
        RECT 4.000 909.520 996.000 910.160 ;
        RECT 4.000 908.120 995.600 909.520 ;
        RECT 4.000 901.360 996.000 908.120 ;
        RECT 4.400 899.960 996.000 901.360 ;
        RECT 4.000 899.320 996.000 899.960 ;
        RECT 4.000 897.920 995.600 899.320 ;
        RECT 4.000 891.160 996.000 897.920 ;
        RECT 4.400 889.760 996.000 891.160 ;
        RECT 4.000 888.440 996.000 889.760 ;
        RECT 4.000 887.040 995.600 888.440 ;
        RECT 4.000 881.640 996.000 887.040 ;
        RECT 4.400 880.240 996.000 881.640 ;
        RECT 4.000 877.560 996.000 880.240 ;
        RECT 4.000 876.160 995.600 877.560 ;
        RECT 4.000 871.440 996.000 876.160 ;
        RECT 4.400 870.040 996.000 871.440 ;
        RECT 4.000 867.360 996.000 870.040 ;
        RECT 4.000 865.960 995.600 867.360 ;
        RECT 4.000 861.240 996.000 865.960 ;
        RECT 4.400 859.840 996.000 861.240 ;
        RECT 4.000 856.480 996.000 859.840 ;
        RECT 4.000 855.080 995.600 856.480 ;
        RECT 4.000 851.040 996.000 855.080 ;
        RECT 4.400 849.640 996.000 851.040 ;
        RECT 4.000 845.600 996.000 849.640 ;
        RECT 4.000 844.200 995.600 845.600 ;
        RECT 4.000 840.840 996.000 844.200 ;
        RECT 4.400 839.440 996.000 840.840 ;
        RECT 4.000 835.400 996.000 839.440 ;
        RECT 4.000 834.000 995.600 835.400 ;
        RECT 4.000 831.320 996.000 834.000 ;
        RECT 4.400 829.920 996.000 831.320 ;
        RECT 4.000 824.520 996.000 829.920 ;
        RECT 4.000 823.120 995.600 824.520 ;
        RECT 4.000 821.120 996.000 823.120 ;
        RECT 4.400 819.720 996.000 821.120 ;
        RECT 4.000 814.320 996.000 819.720 ;
        RECT 4.000 812.920 995.600 814.320 ;
        RECT 4.000 810.920 996.000 812.920 ;
        RECT 4.400 809.520 996.000 810.920 ;
        RECT 4.000 803.440 996.000 809.520 ;
        RECT 4.000 802.040 995.600 803.440 ;
        RECT 4.000 800.720 996.000 802.040 ;
        RECT 4.400 799.320 996.000 800.720 ;
        RECT 4.000 792.560 996.000 799.320 ;
        RECT 4.000 791.160 995.600 792.560 ;
        RECT 4.000 790.520 996.000 791.160 ;
        RECT 4.400 789.120 996.000 790.520 ;
        RECT 4.000 782.360 996.000 789.120 ;
        RECT 4.000 781.000 995.600 782.360 ;
        RECT 4.400 780.960 995.600 781.000 ;
        RECT 4.400 779.600 996.000 780.960 ;
        RECT 4.000 771.480 996.000 779.600 ;
        RECT 4.000 770.800 995.600 771.480 ;
        RECT 4.400 770.080 995.600 770.800 ;
        RECT 4.400 769.400 996.000 770.080 ;
        RECT 4.000 760.600 996.000 769.400 ;
        RECT 4.400 759.200 995.600 760.600 ;
        RECT 4.000 750.400 996.000 759.200 ;
        RECT 4.400 749.000 995.600 750.400 ;
        RECT 4.000 740.200 996.000 749.000 ;
        RECT 4.400 739.520 996.000 740.200 ;
        RECT 4.400 738.800 995.600 739.520 ;
        RECT 4.000 738.120 995.600 738.800 ;
        RECT 4.000 730.000 996.000 738.120 ;
        RECT 4.400 728.640 996.000 730.000 ;
        RECT 4.400 728.600 995.600 728.640 ;
        RECT 4.000 727.240 995.600 728.600 ;
        RECT 4.000 720.480 996.000 727.240 ;
        RECT 4.400 719.080 996.000 720.480 ;
        RECT 4.000 718.440 996.000 719.080 ;
        RECT 4.000 717.040 995.600 718.440 ;
        RECT 4.000 710.280 996.000 717.040 ;
        RECT 4.400 708.880 996.000 710.280 ;
        RECT 4.000 707.560 996.000 708.880 ;
        RECT 4.000 706.160 995.600 707.560 ;
        RECT 4.000 700.080 996.000 706.160 ;
        RECT 4.400 698.680 996.000 700.080 ;
        RECT 4.000 696.680 996.000 698.680 ;
        RECT 4.000 695.280 995.600 696.680 ;
        RECT 4.000 689.880 996.000 695.280 ;
        RECT 4.400 688.480 996.000 689.880 ;
        RECT 4.000 686.480 996.000 688.480 ;
        RECT 4.000 685.080 995.600 686.480 ;
        RECT 4.000 679.680 996.000 685.080 ;
        RECT 4.400 678.280 996.000 679.680 ;
        RECT 4.000 675.600 996.000 678.280 ;
        RECT 4.000 674.200 995.600 675.600 ;
        RECT 4.000 670.160 996.000 674.200 ;
        RECT 4.400 668.760 996.000 670.160 ;
        RECT 4.000 665.400 996.000 668.760 ;
        RECT 4.000 664.000 995.600 665.400 ;
        RECT 4.000 659.960 996.000 664.000 ;
        RECT 4.400 658.560 996.000 659.960 ;
        RECT 4.000 654.520 996.000 658.560 ;
        RECT 4.000 653.120 995.600 654.520 ;
        RECT 4.000 649.760 996.000 653.120 ;
        RECT 4.400 648.360 996.000 649.760 ;
        RECT 4.000 643.640 996.000 648.360 ;
        RECT 4.000 642.240 995.600 643.640 ;
        RECT 4.000 639.560 996.000 642.240 ;
        RECT 4.400 638.160 996.000 639.560 ;
        RECT 4.000 633.440 996.000 638.160 ;
        RECT 4.000 632.040 995.600 633.440 ;
        RECT 4.000 629.360 996.000 632.040 ;
        RECT 4.400 627.960 996.000 629.360 ;
        RECT 4.000 622.560 996.000 627.960 ;
        RECT 4.000 621.160 995.600 622.560 ;
        RECT 4.000 619.840 996.000 621.160 ;
        RECT 4.400 618.440 996.000 619.840 ;
        RECT 4.000 611.680 996.000 618.440 ;
        RECT 4.000 610.280 995.600 611.680 ;
        RECT 4.000 609.640 996.000 610.280 ;
        RECT 4.400 608.240 996.000 609.640 ;
        RECT 4.000 601.480 996.000 608.240 ;
        RECT 4.000 600.080 995.600 601.480 ;
        RECT 4.000 599.440 996.000 600.080 ;
        RECT 4.400 598.040 996.000 599.440 ;
        RECT 4.000 590.600 996.000 598.040 ;
        RECT 4.000 589.240 995.600 590.600 ;
        RECT 4.400 589.200 995.600 589.240 ;
        RECT 4.400 587.840 996.000 589.200 ;
        RECT 4.000 579.720 996.000 587.840 ;
        RECT 4.000 579.040 995.600 579.720 ;
        RECT 4.400 578.320 995.600 579.040 ;
        RECT 4.400 577.640 996.000 578.320 ;
        RECT 4.000 569.520 996.000 577.640 ;
        RECT 4.400 568.120 995.600 569.520 ;
        RECT 4.000 559.320 996.000 568.120 ;
        RECT 4.400 558.640 996.000 559.320 ;
        RECT 4.400 557.920 995.600 558.640 ;
        RECT 4.000 557.240 995.600 557.920 ;
        RECT 4.000 549.120 996.000 557.240 ;
        RECT 4.400 547.760 996.000 549.120 ;
        RECT 4.400 547.720 995.600 547.760 ;
        RECT 4.000 546.360 995.600 547.720 ;
        RECT 4.000 538.920 996.000 546.360 ;
        RECT 4.400 537.560 996.000 538.920 ;
        RECT 4.400 537.520 995.600 537.560 ;
        RECT 4.000 536.160 995.600 537.520 ;
        RECT 4.000 528.720 996.000 536.160 ;
        RECT 4.400 527.320 996.000 528.720 ;
        RECT 4.000 526.680 996.000 527.320 ;
        RECT 4.000 525.280 995.600 526.680 ;
        RECT 4.000 519.200 996.000 525.280 ;
        RECT 4.400 517.800 996.000 519.200 ;
        RECT 4.000 515.800 996.000 517.800 ;
        RECT 4.000 514.400 995.600 515.800 ;
        RECT 4.000 509.000 996.000 514.400 ;
        RECT 4.400 507.600 996.000 509.000 ;
        RECT 4.000 505.600 996.000 507.600 ;
        RECT 4.000 504.200 995.600 505.600 ;
        RECT 4.000 498.800 996.000 504.200 ;
        RECT 4.400 497.400 996.000 498.800 ;
        RECT 4.000 494.720 996.000 497.400 ;
        RECT 4.000 493.320 995.600 494.720 ;
        RECT 4.000 488.600 996.000 493.320 ;
        RECT 4.400 487.200 996.000 488.600 ;
        RECT 4.000 484.520 996.000 487.200 ;
        RECT 4.000 483.120 995.600 484.520 ;
        RECT 4.000 478.400 996.000 483.120 ;
        RECT 4.400 477.000 996.000 478.400 ;
        RECT 4.000 473.640 996.000 477.000 ;
        RECT 4.000 472.240 995.600 473.640 ;
        RECT 4.000 468.880 996.000 472.240 ;
        RECT 4.400 467.480 996.000 468.880 ;
        RECT 4.000 462.760 996.000 467.480 ;
        RECT 4.000 461.360 995.600 462.760 ;
        RECT 4.000 458.680 996.000 461.360 ;
        RECT 4.400 457.280 996.000 458.680 ;
        RECT 4.000 452.560 996.000 457.280 ;
        RECT 4.000 451.160 995.600 452.560 ;
        RECT 4.000 448.480 996.000 451.160 ;
        RECT 4.400 447.080 996.000 448.480 ;
        RECT 4.000 441.680 996.000 447.080 ;
        RECT 4.000 440.280 995.600 441.680 ;
        RECT 4.000 438.280 996.000 440.280 ;
        RECT 4.400 436.880 996.000 438.280 ;
        RECT 4.000 430.800 996.000 436.880 ;
        RECT 4.000 429.400 995.600 430.800 ;
        RECT 4.000 428.080 996.000 429.400 ;
        RECT 4.400 426.680 996.000 428.080 ;
        RECT 4.000 420.600 996.000 426.680 ;
        RECT 4.000 419.200 995.600 420.600 ;
        RECT 4.000 418.560 996.000 419.200 ;
        RECT 4.400 417.160 996.000 418.560 ;
        RECT 4.000 409.720 996.000 417.160 ;
        RECT 4.000 408.360 995.600 409.720 ;
        RECT 4.400 408.320 995.600 408.360 ;
        RECT 4.400 406.960 996.000 408.320 ;
        RECT 4.000 398.840 996.000 406.960 ;
        RECT 4.000 398.160 995.600 398.840 ;
        RECT 4.400 397.440 995.600 398.160 ;
        RECT 4.400 396.760 996.000 397.440 ;
        RECT 4.000 388.640 996.000 396.760 ;
        RECT 4.000 387.960 995.600 388.640 ;
        RECT 4.400 387.240 995.600 387.960 ;
        RECT 4.400 386.560 996.000 387.240 ;
        RECT 4.000 377.760 996.000 386.560 ;
        RECT 4.400 376.360 995.600 377.760 ;
        RECT 4.000 367.560 996.000 376.360 ;
        RECT 4.400 366.880 996.000 367.560 ;
        RECT 4.400 366.160 995.600 366.880 ;
        RECT 4.000 365.480 995.600 366.160 ;
        RECT 4.000 358.040 996.000 365.480 ;
        RECT 4.400 356.680 996.000 358.040 ;
        RECT 4.400 356.640 995.600 356.680 ;
        RECT 4.000 355.280 995.600 356.640 ;
        RECT 4.000 347.840 996.000 355.280 ;
        RECT 4.400 346.440 996.000 347.840 ;
        RECT 4.000 345.800 996.000 346.440 ;
        RECT 4.000 344.400 995.600 345.800 ;
        RECT 4.000 337.640 996.000 344.400 ;
        RECT 4.400 336.240 996.000 337.640 ;
        RECT 4.000 335.600 996.000 336.240 ;
        RECT 4.000 334.200 995.600 335.600 ;
        RECT 4.000 327.440 996.000 334.200 ;
        RECT 4.400 326.040 996.000 327.440 ;
        RECT 4.000 324.720 996.000 326.040 ;
        RECT 4.000 323.320 995.600 324.720 ;
        RECT 4.000 317.240 996.000 323.320 ;
        RECT 4.400 315.840 996.000 317.240 ;
        RECT 4.000 313.840 996.000 315.840 ;
        RECT 4.000 312.440 995.600 313.840 ;
        RECT 4.000 307.720 996.000 312.440 ;
        RECT 4.400 306.320 996.000 307.720 ;
        RECT 4.000 303.640 996.000 306.320 ;
        RECT 4.000 302.240 995.600 303.640 ;
        RECT 4.000 297.520 996.000 302.240 ;
        RECT 4.400 296.120 996.000 297.520 ;
        RECT 4.000 292.760 996.000 296.120 ;
        RECT 4.000 291.360 995.600 292.760 ;
        RECT 4.000 287.320 996.000 291.360 ;
        RECT 4.400 285.920 996.000 287.320 ;
        RECT 4.000 281.880 996.000 285.920 ;
        RECT 4.000 280.480 995.600 281.880 ;
        RECT 4.000 277.120 996.000 280.480 ;
        RECT 4.400 275.720 996.000 277.120 ;
        RECT 4.000 271.680 996.000 275.720 ;
        RECT 4.000 270.280 995.600 271.680 ;
        RECT 4.000 266.920 996.000 270.280 ;
        RECT 4.400 265.520 996.000 266.920 ;
        RECT 4.000 260.800 996.000 265.520 ;
        RECT 4.000 259.400 995.600 260.800 ;
        RECT 4.000 257.400 996.000 259.400 ;
        RECT 4.400 256.000 996.000 257.400 ;
        RECT 4.000 249.920 996.000 256.000 ;
        RECT 4.000 248.520 995.600 249.920 ;
        RECT 4.000 247.200 996.000 248.520 ;
        RECT 4.400 245.800 996.000 247.200 ;
        RECT 4.000 239.720 996.000 245.800 ;
        RECT 4.000 238.320 995.600 239.720 ;
        RECT 4.000 237.000 996.000 238.320 ;
        RECT 4.400 235.600 996.000 237.000 ;
        RECT 4.000 228.840 996.000 235.600 ;
        RECT 4.000 227.440 995.600 228.840 ;
        RECT 4.000 226.800 996.000 227.440 ;
        RECT 4.400 225.400 996.000 226.800 ;
        RECT 4.000 217.960 996.000 225.400 ;
        RECT 4.000 216.600 995.600 217.960 ;
        RECT 4.400 216.560 995.600 216.600 ;
        RECT 4.400 215.200 996.000 216.560 ;
        RECT 4.000 207.760 996.000 215.200 ;
        RECT 4.000 207.080 995.600 207.760 ;
        RECT 4.400 206.360 995.600 207.080 ;
        RECT 4.400 205.680 996.000 206.360 ;
        RECT 4.000 196.880 996.000 205.680 ;
        RECT 4.400 195.480 995.600 196.880 ;
        RECT 4.000 186.680 996.000 195.480 ;
        RECT 4.400 186.000 996.000 186.680 ;
        RECT 4.400 185.280 995.600 186.000 ;
        RECT 4.000 184.600 995.600 185.280 ;
        RECT 4.000 176.480 996.000 184.600 ;
        RECT 4.400 175.800 996.000 176.480 ;
        RECT 4.400 175.080 995.600 175.800 ;
        RECT 4.000 174.400 995.600 175.080 ;
        RECT 4.000 166.280 996.000 174.400 ;
        RECT 4.400 164.920 996.000 166.280 ;
        RECT 4.400 164.880 995.600 164.920 ;
        RECT 4.000 163.520 995.600 164.880 ;
        RECT 4.000 156.760 996.000 163.520 ;
        RECT 4.400 155.360 996.000 156.760 ;
        RECT 4.000 154.720 996.000 155.360 ;
        RECT 4.000 153.320 995.600 154.720 ;
        RECT 4.000 146.560 996.000 153.320 ;
        RECT 4.400 145.160 996.000 146.560 ;
        RECT 4.000 143.840 996.000 145.160 ;
        RECT 4.000 142.440 995.600 143.840 ;
        RECT 4.000 136.360 996.000 142.440 ;
        RECT 4.400 134.960 996.000 136.360 ;
        RECT 4.000 132.960 996.000 134.960 ;
        RECT 4.000 131.560 995.600 132.960 ;
        RECT 4.000 126.160 996.000 131.560 ;
        RECT 4.400 124.760 996.000 126.160 ;
        RECT 4.000 122.760 996.000 124.760 ;
        RECT 4.000 121.360 995.600 122.760 ;
        RECT 4.000 115.960 996.000 121.360 ;
        RECT 4.400 114.560 996.000 115.960 ;
        RECT 4.000 111.880 996.000 114.560 ;
        RECT 4.000 110.480 995.600 111.880 ;
        RECT 4.000 106.440 996.000 110.480 ;
        RECT 4.400 105.040 996.000 106.440 ;
        RECT 4.000 101.000 996.000 105.040 ;
        RECT 4.000 99.600 995.600 101.000 ;
        RECT 4.000 96.240 996.000 99.600 ;
        RECT 4.400 94.840 996.000 96.240 ;
        RECT 4.000 90.800 996.000 94.840 ;
        RECT 4.000 89.400 995.600 90.800 ;
        RECT 4.000 86.040 996.000 89.400 ;
        RECT 4.400 84.640 996.000 86.040 ;
        RECT 4.000 79.920 996.000 84.640 ;
        RECT 4.000 78.520 995.600 79.920 ;
        RECT 4.000 75.840 996.000 78.520 ;
        RECT 4.400 74.440 996.000 75.840 ;
        RECT 4.000 69.040 996.000 74.440 ;
        RECT 4.000 67.640 995.600 69.040 ;
        RECT 4.000 65.640 996.000 67.640 ;
        RECT 4.400 64.240 996.000 65.640 ;
        RECT 4.000 58.840 996.000 64.240 ;
        RECT 4.000 57.440 995.600 58.840 ;
        RECT 4.000 56.120 996.000 57.440 ;
        RECT 4.400 54.720 996.000 56.120 ;
        RECT 4.000 47.960 996.000 54.720 ;
        RECT 4.000 46.560 995.600 47.960 ;
        RECT 4.000 45.920 996.000 46.560 ;
        RECT 4.400 44.520 996.000 45.920 ;
        RECT 4.000 37.080 996.000 44.520 ;
        RECT 4.000 35.720 995.600 37.080 ;
        RECT 4.400 35.680 995.600 35.720 ;
        RECT 4.400 34.320 996.000 35.680 ;
        RECT 4.000 26.880 996.000 34.320 ;
        RECT 4.000 25.520 995.600 26.880 ;
        RECT 4.400 25.480 995.600 25.520 ;
        RECT 4.400 24.120 996.000 25.480 ;
        RECT 4.000 16.000 996.000 24.120 ;
        RECT 4.000 15.320 995.600 16.000 ;
        RECT 4.400 14.600 995.600 15.320 ;
        RECT 4.400 13.920 996.000 14.600 ;
        RECT 4.000 5.800 996.000 13.920 ;
        RECT 4.400 4.935 995.600 5.800 ;
      LAYER met4 ;
        RECT 370.135 26.015 404.640 276.585 ;
        RECT 407.040 26.015 481.440 276.585 ;
        RECT 483.840 26.015 489.145 276.585 ;
  END
END user_proj_example
END LIBRARY

