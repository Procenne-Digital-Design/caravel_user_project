VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 1600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 1596.000 1.750 1600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 1596.000 110.310 1600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 1596.000 120.890 1600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 1596.000 131.930 1600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 1596.000 142.510 1600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 1596.000 153.550 1600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1596.000 164.590 1600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 1596.000 175.170 1600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 1596.000 186.210 1600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1596.000 196.790 1600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 1596.000 207.830 1600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 1596.000 12.330 1600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 1596.000 218.870 1600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 1596.000 229.450 1600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 1596.000 240.490 1600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 1596.000 251.070 1600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 1596.000 262.110 1600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 1596.000 273.150 1600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1596.000 283.730 1600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 1596.000 294.770 1600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 1596.000 305.350 1600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 1596.000 316.390 1600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 1596.000 23.370 1600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 1596.000 327.430 1600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 1596.000 338.010 1600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 1596.000 349.050 1600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 1596.000 360.090 1600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 1596.000 370.670 1600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 1596.000 381.710 1600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 1596.000 392.290 1600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 1596.000 403.330 1600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1596.000 33.950 1600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 1596.000 44.990 1600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 1596.000 56.030 1600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 1596.000 66.610 1600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1596.000 77.650 1600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 1596.000 88.230 1600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 1596.000 99.270 1600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 1596.000 4.970 1600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 1596.000 113.530 1600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 1596.000 124.570 1600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1596.000 135.610 1600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 1596.000 146.190 1600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 1596.000 157.230 1600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1596.000 167.810 1600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 1596.000 178.850 1600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 1596.000 189.890 1600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 1596.000 200.470 1600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 1596.000 211.510 1600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 1596.000 16.010 1600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 1596.000 222.090 1600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 1596.000 233.130 1600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 1596.000 244.170 1600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 1596.000 254.750 1600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 1596.000 265.790 1600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 1596.000 276.830 1600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 1596.000 287.410 1600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 1596.000 298.450 1600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 1596.000 309.030 1600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 1596.000 320.070 1600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 1596.000 27.050 1600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 1596.000 331.110 1600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1596.000 341.690 1600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 1596.000 352.730 1600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 1596.000 363.310 1600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 1596.000 374.350 1600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 1596.000 385.390 1600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 1596.000 395.970 1600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 1596.000 407.010 1600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 1596.000 37.630 1600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1596.000 48.670 1600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 1596.000 59.250 1600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 1596.000 70.290 1600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 1596.000 81.330 1600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 1596.000 91.910 1600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 1596.000 102.950 1600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 1596.000 8.650 1600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 1596.000 117.210 1600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 1596.000 128.250 1600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 1596.000 139.290 1600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 1596.000 149.870 1600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 1596.000 160.910 1600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 1596.000 171.490 1600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 1596.000 182.530 1600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1596.000 193.570 1600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 1596.000 204.150 1600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 1596.000 215.190 1600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1596.000 19.690 1600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1596.000 225.770 1600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 1596.000 236.810 1600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 1596.000 247.850 1600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 1596.000 258.430 1600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 1596.000 269.470 1600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 1596.000 280.050 1600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 1596.000 291.090 1600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 1596.000 302.130 1600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 1596.000 312.710 1600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 1596.000 323.750 1600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 1596.000 30.270 1600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 1596.000 334.330 1600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 1596.000 345.370 1600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 1596.000 356.410 1600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 1596.000 366.990 1600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 1596.000 378.030 1600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 1596.000 388.610 1600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1596.000 399.650 1600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 1596.000 410.690 1600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 1596.000 41.310 1600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 1596.000 52.350 1600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 1596.000 62.930 1600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 1596.000 73.970 1600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 1596.000 84.550 1600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 1596.000 95.590 1600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 1596.000 106.630 1600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1283.200 800.000 1283.800 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.920 4.000 1337.520 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 0.000 752.010 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1358.000 800.000 1358.600 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 1596.000 740.050 1600.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.840 4.000 1418.440 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 278.840 800.000 279.440 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 1596.000 750.630 1600.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 0.000 762.590 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1419.880 800.000 1420.480 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1432.120 800.000 1432.720 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1485.160 4.000 1485.760 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 1596.000 761.670 1600.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1481.760 800.000 1482.360 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1506.920 800.000 1507.520 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 1596.000 775.930 1600.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 1596.000 464.970 1600.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1551.800 4.000 1552.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1531.400 800.000 1532.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 1596.000 783.290 1600.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 0.000 791.110 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 1596.000 790.650 1600.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1568.800 800.000 1569.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 1596.000 798.010 1600.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 303.320 800.000 303.920 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 1596.000 479.230 1600.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 365.200 800.000 365.800 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 1596.000 493.950 1600.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 1596.000 504.530 1600.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 464.480 800.000 465.080 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 489.640 800.000 490.240 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 527.040 800.000 527.640 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.320 4.000 422.920 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 650.800 800.000 651.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 1596.000 551.910 1600.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 92.520 800.000 93.120 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 1596.000 555.130 1600.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 1596.000 562.490 1600.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 762.320 800.000 762.920 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 1596.000 577.210 1600.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 824.200 800.000 824.800 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 1596.000 587.790 1600.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 873.840 800.000 874.440 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 886.760 800.000 887.360 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 911.240 800.000 911.840 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 1596.000 609.410 1600.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 936.400 800.000 937.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 1596.000 616.770 1600.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 948.640 800.000 949.240 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 1596.000 620.450 1600.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 906.480 4.000 907.080 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 1596.000 624.130 1600.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1596.000 631.490 1600.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 1596.000 635.170 1600.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 998.280 800.000 998.880 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1010.520 800.000 1011.120 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 1596.000 645.750 1600.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 1596.000 649.430 1600.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 1596.000 656.790 1600.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 1596.000 660.470 1600.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.120 4.000 1041.720 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.720 4.000 1055.320 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 1596.000 678.410 1600.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1060.160 800.000 1060.760 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1084.640 800.000 1085.240 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 1596.000 685.770 1600.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1097.560 800.000 1098.160 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1109.800 800.000 1110.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1134.280 800.000 1134.880 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 1596.000 696.350 1600.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1229.480 4.000 1230.080 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 229.200 800.000 229.800 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1171.680 800.000 1172.280 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1183.920 800.000 1184.520 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1209.080 800.000 1209.680 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1269.600 4.000 1270.200 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1233.560 800.000 1234.160 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1246.480 800.000 1247.080 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 1596.000 725.330 1600.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1258.720 800.000 1259.320 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 266.600 800.000 267.200 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 18.400 800.000 19.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1295.440 800.000 1296.040 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1308.360 800.000 1308.960 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 1596.000 732.690 1600.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1332.840 800.000 1333.440 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.120 4.000 1364.720 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 1596.000 743.730 1600.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 1596.000 746.950 1600.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 1596.000 754.310 1600.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1407.640 800.000 1408.240 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 1596.000 757.990 1600.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1457.960 4.000 1458.560 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1444.360 800.000 1444.960 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1511.680 4.000 1512.280 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1457.280 800.000 1457.880 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 1596.000 765.350 1600.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 1596.000 769.030 1600.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1525.280 4.000 1525.880 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1538.880 4.000 1539.480 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1565.400 4.000 1566.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1543.640 800.000 1544.240 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 1596.000 786.970 1600.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1581.040 800.000 1581.640 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1593.280 800.000 1593.880 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 340.720 800.000 341.320 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 1596.000 490.270 1600.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 1596.000 497.630 1600.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 1596.000 508.210 1600.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 402.600 800.000 403.200 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 414.840 800.000 415.440 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 1596.000 417.590 1600.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 1596.000 519.250 1600.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 1596.000 522.930 1600.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 501.880 800.000 502.480 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 1596.000 537.190 1600.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 576.680 800.000 577.280 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 601.160 800.000 601.760 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1596.000 544.550 1600.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 1596.000 424.950 1600.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 712.680 800.000 713.280 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 1596.000 558.810 1600.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 1596.000 569.850 1600.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 104.760 800.000 105.360 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1596.000 573.530 1600.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 799.720 800.000 800.320 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 837.120 800.000 837.720 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 849.360 800.000 849.960 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1596.000 584.110 1600.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 1596.000 595.150 1600.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 1596.000 602.510 1600.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 1596.000 439.670 1600.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 4.000 773.120 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 1596.000 446.570 1600.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 1596.000 627.810 1600.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 960.880 800.000 961.480 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 1596.000 638.390 1600.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.000 4.000 1001.600 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 179.560 800.000 180.160 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.920 4.000 1014.520 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1027.520 4.000 1028.120 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1035.000 800.000 1035.600 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1596.000 663.690 1600.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1068.320 4.000 1068.920 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 1596.000 667.370 1600.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 1596.000 671.050 1600.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 1596.000 674.730 1600.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 204.040 800.000 204.640 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 0.000 692.210 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1175.760 4.000 1176.360 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1596.000 689.450 1600.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1147.200 800.000 1147.800 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.280 4.000 1202.880 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 241.440 800.000 242.040 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 1596.000 700.030 1600.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 1596.000 707.390 1600.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1221.320 800.000 1221.920 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 1596.000 714.750 1600.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 1596.000 718.430 1600.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.720 4.000 1310.320 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1270.960 800.000 1271.560 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 1596.000 461.290 1600.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1323.320 4.000 1323.920 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 1596.000 729.010 1600.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1320.600 800.000 1321.200 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1350.520 4.000 1351.120 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1345.080 800.000 1345.680 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1370.240 800.000 1370.840 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 1596.000 736.370 1600.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1382.480 800.000 1383.080 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1394.720 800.000 1395.320 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.760 4.000 1431.360 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1444.360 4.000 1444.960 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1471.560 4.000 1472.160 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.080 4.000 1498.680 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1469.520 800.000 1470.120 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1494.000 800.000 1494.600 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 1596.000 772.710 1600.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1519.160 800.000 1519.760 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 1596.000 468.650 1600.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1596.000 779.610 1600.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1556.560 800.000 1557.160 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1579.000 4.000 1579.600 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 1596.000 794.330 1600.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1592.600 4.000 1593.200 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 1596.000 475.550 1600.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 1596.000 482.910 1600.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 378.120 800.000 378.720 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 1596.000 511.890 1600.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 1596.000 421.270 1600.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 477.400 800.000 478.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 1596.000 529.830 1600.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 539.280 800.000 539.880 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 613.400 800.000 614.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 626.320 800.000 626.920 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 1596.000 548.230 1600.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 675.280 800.000 675.880 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.160 4.000 584.760 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 724.920 800.000 725.520 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 737.840 800.000 738.440 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 750.080 800.000 750.680 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 1596.000 566.170 1600.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 774.560 800.000 775.160 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 787.480 800.000 788.080 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 811.960 800.000 812.560 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 1596.000 580.890 1600.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 861.600 800.000 862.200 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 1596.000 591.470 1600.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 1596.000 598.830 1600.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 1596.000 442.890 1600.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 899.000 800.000 899.600 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 1596.000 606.190 1600.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 923.480 800.000 924.080 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 1596.000 613.090 1600.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 4.000 853.360 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 142.160 800.000 142.760 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.680 4.000 934.280 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.280 4.000 947.880 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 973.120 800.000 973.720 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 985.360 800.000 985.960 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.800 4.000 974.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 1596.000 642.070 1600.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 1596.000 653.110 1600.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1022.760 800.000 1023.360 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1047.920 800.000 1048.520 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 4.000 1135.560 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1148.560 4.000 1149.160 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 216.960 800.000 217.560 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1072.400 800.000 1073.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 1596.000 682.090 1600.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1189.360 4.000 1189.960 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1122.040 800.000 1122.640 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1596.000 692.670 1600.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.880 4.000 1216.480 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1159.440 800.000 1160.040 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1256.000 4.000 1256.600 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1196.840 800.000 1197.440 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 1596.000 703.710 1600.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 1596.000 711.070 1600.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1283.200 4.000 1283.800 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1296.800 4.000 1297.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1596.000 721.650 1600.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END la_oenb[9]
  PIN sram_addr_a[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 30.640 800.000 31.240 ;
    END
  END sram_addr_a[0]
  PIN sram_addr_a[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END sram_addr_a[1]
  PIN sram_addr_a[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END sram_addr_a[2]
  PIN sram_addr_a[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 1596.000 432.310 1600.000 ;
    END
  END sram_addr_a[3]
  PIN sram_addr_a[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 129.920 800.000 130.520 ;
    END
  END sram_addr_a[4]
  PIN sram_addr_a[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END sram_addr_a[5]
  PIN sram_addr_a[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END sram_addr_a[6]
  PIN sram_addr_a[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END sram_addr_a[7]
  PIN sram_addr_a[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END sram_addr_a[8]
  PIN sram_addr_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 42.880 800.000 43.480 ;
    END
  END sram_addr_b[0]
  PIN sram_addr_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END sram_addr_b[1]
  PIN sram_addr_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END sram_addr_b[2]
  PIN sram_addr_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 1596.000 435.990 1600.000 ;
    END
  END sram_addr_b[3]
  PIN sram_addr_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END sram_addr_b[4]
  PIN sram_addr_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 154.400 800.000 155.000 ;
    END
  END sram_addr_b[5]
  PIN sram_addr_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 1596.000 450.250 1600.000 ;
    END
  END sram_addr_b[6]
  PIN sram_addr_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END sram_addr_b[7]
  PIN sram_addr_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 1596.000 457.610 1600.000 ;
    END
  END sram_addr_b[8]
  PIN sram_csb_a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 6.160 800.000 6.760 ;
    END
  END sram_csb_a
  PIN sram_csb_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END sram_csb_b
  PIN sram_din_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END sram_din_b[0]
  PIN sram_din_b[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END sram_din_b[10]
  PIN sram_din_b[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END sram_din_b[11]
  PIN sram_din_b[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 316.240 800.000 316.840 ;
    END
  END sram_din_b[12]
  PIN sram_din_b[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 1596.000 486.590 1600.000 ;
    END
  END sram_din_b[13]
  PIN sram_din_b[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END sram_din_b[14]
  PIN sram_din_b[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END sram_din_b[15]
  PIN sram_din_b[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END sram_din_b[16]
  PIN sram_din_b[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END sram_din_b[17]
  PIN sram_din_b[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END sram_din_b[18]
  PIN sram_din_b[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END sram_din_b[19]
  PIN sram_din_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 55.120 800.000 55.720 ;
    END
  END sram_din_b[1]
  PIN sram_din_b[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 440.000 800.000 440.600 ;
    END
  END sram_din_b[20]
  PIN sram_din_b[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 452.240 800.000 452.840 ;
    END
  END sram_din_b[21]
  PIN sram_din_b[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 1596.000 526.150 1600.000 ;
    END
  END sram_din_b[22]
  PIN sram_din_b[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 514.120 800.000 514.720 ;
    END
  END sram_din_b[23]
  PIN sram_din_b[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 551.520 800.000 552.120 ;
    END
  END sram_din_b[24]
  PIN sram_din_b[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 588.920 800.000 589.520 ;
    END
  END sram_din_b[25]
  PIN sram_din_b[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END sram_din_b[26]
  PIN sram_din_b[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END sram_din_b[27]
  PIN sram_din_b[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END sram_din_b[28]
  PIN sram_din_b[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END sram_din_b[29]
  PIN sram_din_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END sram_din_b[2]
  PIN sram_din_b[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 688.200 800.000 688.800 ;
    END
  END sram_din_b[30]
  PIN sram_din_b[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END sram_din_b[31]
  PIN sram_din_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END sram_din_b[3]
  PIN sram_din_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END sram_din_b[4]
  PIN sram_din_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 167.320 800.000 167.920 ;
    END
  END sram_din_b[5]
  PIN sram_din_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 191.800 800.000 192.400 ;
    END
  END sram_din_b[6]
  PIN sram_din_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 1596.000 453.930 1600.000 ;
    END
  END sram_din_b[7]
  PIN sram_din_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END sram_din_b[8]
  PIN sram_din_b[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END sram_din_b[9]
  PIN sram_dout_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END sram_dout_a[0]
  PIN sram_dout_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 291.080 800.000 291.680 ;
    END
  END sram_dout_a[10]
  PIN sram_dout_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 1596.000 471.870 1600.000 ;
    END
  END sram_dout_a[11]
  PIN sram_dout_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 328.480 800.000 329.080 ;
    END
  END sram_dout_a[12]
  PIN sram_dout_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 352.960 800.000 353.560 ;
    END
  END sram_dout_a[13]
  PIN sram_dout_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END sram_dout_a[14]
  PIN sram_dout_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END sram_dout_a[15]
  PIN sram_dout_a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 1596.000 500.850 1600.000 ;
    END
  END sram_dout_a[16]
  PIN sram_dout_a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 390.360 800.000 390.960 ;
    END
  END sram_dout_a[17]
  PIN sram_dout_a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 1596.000 515.570 1600.000 ;
    END
  END sram_dout_a[18]
  PIN sram_dout_a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 427.760 800.000 428.360 ;
    END
  END sram_dout_a[19]
  PIN sram_dout_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 68.040 800.000 68.640 ;
    END
  END sram_dout_a[1]
  PIN sram_dout_a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END sram_dout_a[20]
  PIN sram_dout_a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END sram_dout_a[21]
  PIN sram_dout_a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END sram_dout_a[22]
  PIN sram_dout_a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 1596.000 533.510 1600.000 ;
    END
  END sram_dout_a[23]
  PIN sram_dout_a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 563.760 800.000 564.360 ;
    END
  END sram_dout_a[24]
  PIN sram_dout_a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END sram_dout_a[25]
  PIN sram_dout_a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 1596.000 540.870 1600.000 ;
    END
  END sram_dout_a[26]
  PIN sram_dout_a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 638.560 800.000 639.160 ;
    END
  END sram_dout_a[27]
  PIN sram_dout_a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 663.040 800.000 663.640 ;
    END
  END sram_dout_a[28]
  PIN sram_dout_a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END sram_dout_a[29]
  PIN sram_dout_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1596.000 428.630 1600.000 ;
    END
  END sram_dout_a[2]
  PIN sram_dout_a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 700.440 800.000 701.040 ;
    END
  END sram_dout_a[30]
  PIN sram_dout_a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END sram_dout_a[31]
  PIN sram_dout_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END sram_dout_a[3]
  PIN sram_dout_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END sram_dout_a[4]
  PIN sram_dout_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END sram_dout_a[5]
  PIN sram_dout_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END sram_dout_a[6]
  PIN sram_dout_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END sram_dout_a[7]
  PIN sram_dout_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 253.680 800.000 254.280 ;
    END
  END sram_dout_a[8]
  PIN sram_dout_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END sram_dout_a[9]
  PIN sram_mask_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 1596.000 414.370 1600.000 ;
    END
  END sram_mask_b[0]
  PIN sram_mask_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 80.280 800.000 80.880 ;
    END
  END sram_mask_b[1]
  PIN sram_mask_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END sram_mask_b[2]
  PIN sram_mask_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 117.680 800.000 118.280 ;
    END
  END sram_mask_b[3]
  PIN sram_web_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END sram_web_b
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1588.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1588.720 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 1588.565 ;
      LAYER met1 ;
        RECT 0.070 5.480 798.030 1588.720 ;
      LAYER met2 ;
        RECT 0.100 1595.720 1.190 1596.370 ;
        RECT 2.030 1595.720 4.410 1596.370 ;
        RECT 5.250 1595.720 8.090 1596.370 ;
        RECT 8.930 1595.720 11.770 1596.370 ;
        RECT 12.610 1595.720 15.450 1596.370 ;
        RECT 16.290 1595.720 19.130 1596.370 ;
        RECT 19.970 1595.720 22.810 1596.370 ;
        RECT 23.650 1595.720 26.490 1596.370 ;
        RECT 27.330 1595.720 29.710 1596.370 ;
        RECT 30.550 1595.720 33.390 1596.370 ;
        RECT 34.230 1595.720 37.070 1596.370 ;
        RECT 37.910 1595.720 40.750 1596.370 ;
        RECT 41.590 1595.720 44.430 1596.370 ;
        RECT 45.270 1595.720 48.110 1596.370 ;
        RECT 48.950 1595.720 51.790 1596.370 ;
        RECT 52.630 1595.720 55.470 1596.370 ;
        RECT 56.310 1595.720 58.690 1596.370 ;
        RECT 59.530 1595.720 62.370 1596.370 ;
        RECT 63.210 1595.720 66.050 1596.370 ;
        RECT 66.890 1595.720 69.730 1596.370 ;
        RECT 70.570 1595.720 73.410 1596.370 ;
        RECT 74.250 1595.720 77.090 1596.370 ;
        RECT 77.930 1595.720 80.770 1596.370 ;
        RECT 81.610 1595.720 83.990 1596.370 ;
        RECT 84.830 1595.720 87.670 1596.370 ;
        RECT 88.510 1595.720 91.350 1596.370 ;
        RECT 92.190 1595.720 95.030 1596.370 ;
        RECT 95.870 1595.720 98.710 1596.370 ;
        RECT 99.550 1595.720 102.390 1596.370 ;
        RECT 103.230 1595.720 106.070 1596.370 ;
        RECT 106.910 1595.720 109.750 1596.370 ;
        RECT 110.590 1595.720 112.970 1596.370 ;
        RECT 113.810 1595.720 116.650 1596.370 ;
        RECT 117.490 1595.720 120.330 1596.370 ;
        RECT 121.170 1595.720 124.010 1596.370 ;
        RECT 124.850 1595.720 127.690 1596.370 ;
        RECT 128.530 1595.720 131.370 1596.370 ;
        RECT 132.210 1595.720 135.050 1596.370 ;
        RECT 135.890 1595.720 138.730 1596.370 ;
        RECT 139.570 1595.720 141.950 1596.370 ;
        RECT 142.790 1595.720 145.630 1596.370 ;
        RECT 146.470 1595.720 149.310 1596.370 ;
        RECT 150.150 1595.720 152.990 1596.370 ;
        RECT 153.830 1595.720 156.670 1596.370 ;
        RECT 157.510 1595.720 160.350 1596.370 ;
        RECT 161.190 1595.720 164.030 1596.370 ;
        RECT 164.870 1595.720 167.250 1596.370 ;
        RECT 168.090 1595.720 170.930 1596.370 ;
        RECT 171.770 1595.720 174.610 1596.370 ;
        RECT 175.450 1595.720 178.290 1596.370 ;
        RECT 179.130 1595.720 181.970 1596.370 ;
        RECT 182.810 1595.720 185.650 1596.370 ;
        RECT 186.490 1595.720 189.330 1596.370 ;
        RECT 190.170 1595.720 193.010 1596.370 ;
        RECT 193.850 1595.720 196.230 1596.370 ;
        RECT 197.070 1595.720 199.910 1596.370 ;
        RECT 200.750 1595.720 203.590 1596.370 ;
        RECT 204.430 1595.720 207.270 1596.370 ;
        RECT 208.110 1595.720 210.950 1596.370 ;
        RECT 211.790 1595.720 214.630 1596.370 ;
        RECT 215.470 1595.720 218.310 1596.370 ;
        RECT 219.150 1595.720 221.530 1596.370 ;
        RECT 222.370 1595.720 225.210 1596.370 ;
        RECT 226.050 1595.720 228.890 1596.370 ;
        RECT 229.730 1595.720 232.570 1596.370 ;
        RECT 233.410 1595.720 236.250 1596.370 ;
        RECT 237.090 1595.720 239.930 1596.370 ;
        RECT 240.770 1595.720 243.610 1596.370 ;
        RECT 244.450 1595.720 247.290 1596.370 ;
        RECT 248.130 1595.720 250.510 1596.370 ;
        RECT 251.350 1595.720 254.190 1596.370 ;
        RECT 255.030 1595.720 257.870 1596.370 ;
        RECT 258.710 1595.720 261.550 1596.370 ;
        RECT 262.390 1595.720 265.230 1596.370 ;
        RECT 266.070 1595.720 268.910 1596.370 ;
        RECT 269.750 1595.720 272.590 1596.370 ;
        RECT 273.430 1595.720 276.270 1596.370 ;
        RECT 277.110 1595.720 279.490 1596.370 ;
        RECT 280.330 1595.720 283.170 1596.370 ;
        RECT 284.010 1595.720 286.850 1596.370 ;
        RECT 287.690 1595.720 290.530 1596.370 ;
        RECT 291.370 1595.720 294.210 1596.370 ;
        RECT 295.050 1595.720 297.890 1596.370 ;
        RECT 298.730 1595.720 301.570 1596.370 ;
        RECT 302.410 1595.720 304.790 1596.370 ;
        RECT 305.630 1595.720 308.470 1596.370 ;
        RECT 309.310 1595.720 312.150 1596.370 ;
        RECT 312.990 1595.720 315.830 1596.370 ;
        RECT 316.670 1595.720 319.510 1596.370 ;
        RECT 320.350 1595.720 323.190 1596.370 ;
        RECT 324.030 1595.720 326.870 1596.370 ;
        RECT 327.710 1595.720 330.550 1596.370 ;
        RECT 331.390 1595.720 333.770 1596.370 ;
        RECT 334.610 1595.720 337.450 1596.370 ;
        RECT 338.290 1595.720 341.130 1596.370 ;
        RECT 341.970 1595.720 344.810 1596.370 ;
        RECT 345.650 1595.720 348.490 1596.370 ;
        RECT 349.330 1595.720 352.170 1596.370 ;
        RECT 353.010 1595.720 355.850 1596.370 ;
        RECT 356.690 1595.720 359.530 1596.370 ;
        RECT 360.370 1595.720 362.750 1596.370 ;
        RECT 363.590 1595.720 366.430 1596.370 ;
        RECT 367.270 1595.720 370.110 1596.370 ;
        RECT 370.950 1595.720 373.790 1596.370 ;
        RECT 374.630 1595.720 377.470 1596.370 ;
        RECT 378.310 1595.720 381.150 1596.370 ;
        RECT 381.990 1595.720 384.830 1596.370 ;
        RECT 385.670 1595.720 388.050 1596.370 ;
        RECT 388.890 1595.720 391.730 1596.370 ;
        RECT 392.570 1595.720 395.410 1596.370 ;
        RECT 396.250 1595.720 399.090 1596.370 ;
        RECT 399.930 1595.720 402.770 1596.370 ;
        RECT 403.610 1595.720 406.450 1596.370 ;
        RECT 407.290 1595.720 410.130 1596.370 ;
        RECT 410.970 1595.720 413.810 1596.370 ;
        RECT 414.650 1595.720 417.030 1596.370 ;
        RECT 417.870 1595.720 420.710 1596.370 ;
        RECT 421.550 1595.720 424.390 1596.370 ;
        RECT 425.230 1595.720 428.070 1596.370 ;
        RECT 428.910 1595.720 431.750 1596.370 ;
        RECT 432.590 1595.720 435.430 1596.370 ;
        RECT 436.270 1595.720 439.110 1596.370 ;
        RECT 439.950 1595.720 442.330 1596.370 ;
        RECT 443.170 1595.720 446.010 1596.370 ;
        RECT 446.850 1595.720 449.690 1596.370 ;
        RECT 450.530 1595.720 453.370 1596.370 ;
        RECT 454.210 1595.720 457.050 1596.370 ;
        RECT 457.890 1595.720 460.730 1596.370 ;
        RECT 461.570 1595.720 464.410 1596.370 ;
        RECT 465.250 1595.720 468.090 1596.370 ;
        RECT 468.930 1595.720 471.310 1596.370 ;
        RECT 472.150 1595.720 474.990 1596.370 ;
        RECT 475.830 1595.720 478.670 1596.370 ;
        RECT 479.510 1595.720 482.350 1596.370 ;
        RECT 483.190 1595.720 486.030 1596.370 ;
        RECT 486.870 1595.720 489.710 1596.370 ;
        RECT 490.550 1595.720 493.390 1596.370 ;
        RECT 494.230 1595.720 497.070 1596.370 ;
        RECT 497.910 1595.720 500.290 1596.370 ;
        RECT 501.130 1595.720 503.970 1596.370 ;
        RECT 504.810 1595.720 507.650 1596.370 ;
        RECT 508.490 1595.720 511.330 1596.370 ;
        RECT 512.170 1595.720 515.010 1596.370 ;
        RECT 515.850 1595.720 518.690 1596.370 ;
        RECT 519.530 1595.720 522.370 1596.370 ;
        RECT 523.210 1595.720 525.590 1596.370 ;
        RECT 526.430 1595.720 529.270 1596.370 ;
        RECT 530.110 1595.720 532.950 1596.370 ;
        RECT 533.790 1595.720 536.630 1596.370 ;
        RECT 537.470 1595.720 540.310 1596.370 ;
        RECT 541.150 1595.720 543.990 1596.370 ;
        RECT 544.830 1595.720 547.670 1596.370 ;
        RECT 548.510 1595.720 551.350 1596.370 ;
        RECT 552.190 1595.720 554.570 1596.370 ;
        RECT 555.410 1595.720 558.250 1596.370 ;
        RECT 559.090 1595.720 561.930 1596.370 ;
        RECT 562.770 1595.720 565.610 1596.370 ;
        RECT 566.450 1595.720 569.290 1596.370 ;
        RECT 570.130 1595.720 572.970 1596.370 ;
        RECT 573.810 1595.720 576.650 1596.370 ;
        RECT 577.490 1595.720 580.330 1596.370 ;
        RECT 581.170 1595.720 583.550 1596.370 ;
        RECT 584.390 1595.720 587.230 1596.370 ;
        RECT 588.070 1595.720 590.910 1596.370 ;
        RECT 591.750 1595.720 594.590 1596.370 ;
        RECT 595.430 1595.720 598.270 1596.370 ;
        RECT 599.110 1595.720 601.950 1596.370 ;
        RECT 602.790 1595.720 605.630 1596.370 ;
        RECT 606.470 1595.720 608.850 1596.370 ;
        RECT 609.690 1595.720 612.530 1596.370 ;
        RECT 613.370 1595.720 616.210 1596.370 ;
        RECT 617.050 1595.720 619.890 1596.370 ;
        RECT 620.730 1595.720 623.570 1596.370 ;
        RECT 624.410 1595.720 627.250 1596.370 ;
        RECT 628.090 1595.720 630.930 1596.370 ;
        RECT 631.770 1595.720 634.610 1596.370 ;
        RECT 635.450 1595.720 637.830 1596.370 ;
        RECT 638.670 1595.720 641.510 1596.370 ;
        RECT 642.350 1595.720 645.190 1596.370 ;
        RECT 646.030 1595.720 648.870 1596.370 ;
        RECT 649.710 1595.720 652.550 1596.370 ;
        RECT 653.390 1595.720 656.230 1596.370 ;
        RECT 657.070 1595.720 659.910 1596.370 ;
        RECT 660.750 1595.720 663.130 1596.370 ;
        RECT 663.970 1595.720 666.810 1596.370 ;
        RECT 667.650 1595.720 670.490 1596.370 ;
        RECT 671.330 1595.720 674.170 1596.370 ;
        RECT 675.010 1595.720 677.850 1596.370 ;
        RECT 678.690 1595.720 681.530 1596.370 ;
        RECT 682.370 1595.720 685.210 1596.370 ;
        RECT 686.050 1595.720 688.890 1596.370 ;
        RECT 689.730 1595.720 692.110 1596.370 ;
        RECT 692.950 1595.720 695.790 1596.370 ;
        RECT 696.630 1595.720 699.470 1596.370 ;
        RECT 700.310 1595.720 703.150 1596.370 ;
        RECT 703.990 1595.720 706.830 1596.370 ;
        RECT 707.670 1595.720 710.510 1596.370 ;
        RECT 711.350 1595.720 714.190 1596.370 ;
        RECT 715.030 1595.720 717.870 1596.370 ;
        RECT 718.710 1595.720 721.090 1596.370 ;
        RECT 721.930 1595.720 724.770 1596.370 ;
        RECT 725.610 1595.720 728.450 1596.370 ;
        RECT 729.290 1595.720 732.130 1596.370 ;
        RECT 732.970 1595.720 735.810 1596.370 ;
        RECT 736.650 1595.720 739.490 1596.370 ;
        RECT 740.330 1595.720 743.170 1596.370 ;
        RECT 744.010 1595.720 746.390 1596.370 ;
        RECT 747.230 1595.720 750.070 1596.370 ;
        RECT 750.910 1595.720 753.750 1596.370 ;
        RECT 754.590 1595.720 757.430 1596.370 ;
        RECT 758.270 1595.720 761.110 1596.370 ;
        RECT 761.950 1595.720 764.790 1596.370 ;
        RECT 765.630 1595.720 768.470 1596.370 ;
        RECT 769.310 1595.720 772.150 1596.370 ;
        RECT 772.990 1595.720 775.370 1596.370 ;
        RECT 776.210 1595.720 779.050 1596.370 ;
        RECT 779.890 1595.720 782.730 1596.370 ;
        RECT 783.570 1595.720 786.410 1596.370 ;
        RECT 787.250 1595.720 790.090 1596.370 ;
        RECT 790.930 1595.720 793.770 1596.370 ;
        RECT 794.610 1595.720 797.450 1596.370 ;
        RECT 0.100 4.280 798.000 1595.720 ;
        RECT 0.100 3.670 1.190 4.280 ;
        RECT 2.030 3.670 4.410 4.280 ;
        RECT 5.250 3.670 8.090 4.280 ;
        RECT 8.930 3.670 11.310 4.280 ;
        RECT 12.150 3.670 14.990 4.280 ;
        RECT 15.830 3.670 18.670 4.280 ;
        RECT 19.510 3.670 21.890 4.280 ;
        RECT 22.730 3.670 25.570 4.280 ;
        RECT 26.410 3.670 29.250 4.280 ;
        RECT 30.090 3.670 32.470 4.280 ;
        RECT 33.310 3.670 36.150 4.280 ;
        RECT 36.990 3.670 39.830 4.280 ;
        RECT 40.670 3.670 43.050 4.280 ;
        RECT 43.890 3.670 46.730 4.280 ;
        RECT 47.570 3.670 50.410 4.280 ;
        RECT 51.250 3.670 53.630 4.280 ;
        RECT 54.470 3.670 57.310 4.280 ;
        RECT 58.150 3.670 60.990 4.280 ;
        RECT 61.830 3.670 64.210 4.280 ;
        RECT 65.050 3.670 67.890 4.280 ;
        RECT 68.730 3.670 71.570 4.280 ;
        RECT 72.410 3.670 74.790 4.280 ;
        RECT 75.630 3.670 78.470 4.280 ;
        RECT 79.310 3.670 82.150 4.280 ;
        RECT 82.990 3.670 85.370 4.280 ;
        RECT 86.210 3.670 89.050 4.280 ;
        RECT 89.890 3.670 92.730 4.280 ;
        RECT 93.570 3.670 95.950 4.280 ;
        RECT 96.790 3.670 99.630 4.280 ;
        RECT 100.470 3.670 103.310 4.280 ;
        RECT 104.150 3.670 106.530 4.280 ;
        RECT 107.370 3.670 110.210 4.280 ;
        RECT 111.050 3.670 113.890 4.280 ;
        RECT 114.730 3.670 117.110 4.280 ;
        RECT 117.950 3.670 120.790 4.280 ;
        RECT 121.630 3.670 124.470 4.280 ;
        RECT 125.310 3.670 127.690 4.280 ;
        RECT 128.530 3.670 131.370 4.280 ;
        RECT 132.210 3.670 135.050 4.280 ;
        RECT 135.890 3.670 138.270 4.280 ;
        RECT 139.110 3.670 141.950 4.280 ;
        RECT 142.790 3.670 145.630 4.280 ;
        RECT 146.470 3.670 148.850 4.280 ;
        RECT 149.690 3.670 152.530 4.280 ;
        RECT 153.370 3.670 156.210 4.280 ;
        RECT 157.050 3.670 159.430 4.280 ;
        RECT 160.270 3.670 163.110 4.280 ;
        RECT 163.950 3.670 166.790 4.280 ;
        RECT 167.630 3.670 170.010 4.280 ;
        RECT 170.850 3.670 173.690 4.280 ;
        RECT 174.530 3.670 177.370 4.280 ;
        RECT 178.210 3.670 180.590 4.280 ;
        RECT 181.430 3.670 184.270 4.280 ;
        RECT 185.110 3.670 187.950 4.280 ;
        RECT 188.790 3.670 191.170 4.280 ;
        RECT 192.010 3.670 194.850 4.280 ;
        RECT 195.690 3.670 198.530 4.280 ;
        RECT 199.370 3.670 201.750 4.280 ;
        RECT 202.590 3.670 205.430 4.280 ;
        RECT 206.270 3.670 208.650 4.280 ;
        RECT 209.490 3.670 212.330 4.280 ;
        RECT 213.170 3.670 216.010 4.280 ;
        RECT 216.850 3.670 219.230 4.280 ;
        RECT 220.070 3.670 222.910 4.280 ;
        RECT 223.750 3.670 226.590 4.280 ;
        RECT 227.430 3.670 229.810 4.280 ;
        RECT 230.650 3.670 233.490 4.280 ;
        RECT 234.330 3.670 237.170 4.280 ;
        RECT 238.010 3.670 240.390 4.280 ;
        RECT 241.230 3.670 244.070 4.280 ;
        RECT 244.910 3.670 247.750 4.280 ;
        RECT 248.590 3.670 250.970 4.280 ;
        RECT 251.810 3.670 254.650 4.280 ;
        RECT 255.490 3.670 258.330 4.280 ;
        RECT 259.170 3.670 261.550 4.280 ;
        RECT 262.390 3.670 265.230 4.280 ;
        RECT 266.070 3.670 268.910 4.280 ;
        RECT 269.750 3.670 272.130 4.280 ;
        RECT 272.970 3.670 275.810 4.280 ;
        RECT 276.650 3.670 279.490 4.280 ;
        RECT 280.330 3.670 282.710 4.280 ;
        RECT 283.550 3.670 286.390 4.280 ;
        RECT 287.230 3.670 290.070 4.280 ;
        RECT 290.910 3.670 293.290 4.280 ;
        RECT 294.130 3.670 296.970 4.280 ;
        RECT 297.810 3.670 300.650 4.280 ;
        RECT 301.490 3.670 303.870 4.280 ;
        RECT 304.710 3.670 307.550 4.280 ;
        RECT 308.390 3.670 311.230 4.280 ;
        RECT 312.070 3.670 314.450 4.280 ;
        RECT 315.290 3.670 318.130 4.280 ;
        RECT 318.970 3.670 321.810 4.280 ;
        RECT 322.650 3.670 325.030 4.280 ;
        RECT 325.870 3.670 328.710 4.280 ;
        RECT 329.550 3.670 332.390 4.280 ;
        RECT 333.230 3.670 335.610 4.280 ;
        RECT 336.450 3.670 339.290 4.280 ;
        RECT 340.130 3.670 342.970 4.280 ;
        RECT 343.810 3.670 346.190 4.280 ;
        RECT 347.030 3.670 349.870 4.280 ;
        RECT 350.710 3.670 353.550 4.280 ;
        RECT 354.390 3.670 356.770 4.280 ;
        RECT 357.610 3.670 360.450 4.280 ;
        RECT 361.290 3.670 364.130 4.280 ;
        RECT 364.970 3.670 367.350 4.280 ;
        RECT 368.190 3.670 371.030 4.280 ;
        RECT 371.870 3.670 374.710 4.280 ;
        RECT 375.550 3.670 377.930 4.280 ;
        RECT 378.770 3.670 381.610 4.280 ;
        RECT 382.450 3.670 385.290 4.280 ;
        RECT 386.130 3.670 388.510 4.280 ;
        RECT 389.350 3.670 392.190 4.280 ;
        RECT 393.030 3.670 395.870 4.280 ;
        RECT 396.710 3.670 399.090 4.280 ;
        RECT 399.930 3.670 402.770 4.280 ;
        RECT 403.610 3.670 405.990 4.280 ;
        RECT 406.830 3.670 409.670 4.280 ;
        RECT 410.510 3.670 413.350 4.280 ;
        RECT 414.190 3.670 416.570 4.280 ;
        RECT 417.410 3.670 420.250 4.280 ;
        RECT 421.090 3.670 423.930 4.280 ;
        RECT 424.770 3.670 427.150 4.280 ;
        RECT 427.990 3.670 430.830 4.280 ;
        RECT 431.670 3.670 434.510 4.280 ;
        RECT 435.350 3.670 437.730 4.280 ;
        RECT 438.570 3.670 441.410 4.280 ;
        RECT 442.250 3.670 445.090 4.280 ;
        RECT 445.930 3.670 448.310 4.280 ;
        RECT 449.150 3.670 451.990 4.280 ;
        RECT 452.830 3.670 455.670 4.280 ;
        RECT 456.510 3.670 458.890 4.280 ;
        RECT 459.730 3.670 462.570 4.280 ;
        RECT 463.410 3.670 466.250 4.280 ;
        RECT 467.090 3.670 469.470 4.280 ;
        RECT 470.310 3.670 473.150 4.280 ;
        RECT 473.990 3.670 476.830 4.280 ;
        RECT 477.670 3.670 480.050 4.280 ;
        RECT 480.890 3.670 483.730 4.280 ;
        RECT 484.570 3.670 487.410 4.280 ;
        RECT 488.250 3.670 490.630 4.280 ;
        RECT 491.470 3.670 494.310 4.280 ;
        RECT 495.150 3.670 497.990 4.280 ;
        RECT 498.830 3.670 501.210 4.280 ;
        RECT 502.050 3.670 504.890 4.280 ;
        RECT 505.730 3.670 508.570 4.280 ;
        RECT 509.410 3.670 511.790 4.280 ;
        RECT 512.630 3.670 515.470 4.280 ;
        RECT 516.310 3.670 519.150 4.280 ;
        RECT 519.990 3.670 522.370 4.280 ;
        RECT 523.210 3.670 526.050 4.280 ;
        RECT 526.890 3.670 529.730 4.280 ;
        RECT 530.570 3.670 532.950 4.280 ;
        RECT 533.790 3.670 536.630 4.280 ;
        RECT 537.470 3.670 540.310 4.280 ;
        RECT 541.150 3.670 543.530 4.280 ;
        RECT 544.370 3.670 547.210 4.280 ;
        RECT 548.050 3.670 550.890 4.280 ;
        RECT 551.730 3.670 554.110 4.280 ;
        RECT 554.950 3.670 557.790 4.280 ;
        RECT 558.630 3.670 561.470 4.280 ;
        RECT 562.310 3.670 564.690 4.280 ;
        RECT 565.530 3.670 568.370 4.280 ;
        RECT 569.210 3.670 572.050 4.280 ;
        RECT 572.890 3.670 575.270 4.280 ;
        RECT 576.110 3.670 578.950 4.280 ;
        RECT 579.790 3.670 582.630 4.280 ;
        RECT 583.470 3.670 585.850 4.280 ;
        RECT 586.690 3.670 589.530 4.280 ;
        RECT 590.370 3.670 593.210 4.280 ;
        RECT 594.050 3.670 596.430 4.280 ;
        RECT 597.270 3.670 600.110 4.280 ;
        RECT 600.950 3.670 603.330 4.280 ;
        RECT 604.170 3.670 607.010 4.280 ;
        RECT 607.850 3.670 610.690 4.280 ;
        RECT 611.530 3.670 613.910 4.280 ;
        RECT 614.750 3.670 617.590 4.280 ;
        RECT 618.430 3.670 621.270 4.280 ;
        RECT 622.110 3.670 624.490 4.280 ;
        RECT 625.330 3.670 628.170 4.280 ;
        RECT 629.010 3.670 631.850 4.280 ;
        RECT 632.690 3.670 635.070 4.280 ;
        RECT 635.910 3.670 638.750 4.280 ;
        RECT 639.590 3.670 642.430 4.280 ;
        RECT 643.270 3.670 645.650 4.280 ;
        RECT 646.490 3.670 649.330 4.280 ;
        RECT 650.170 3.670 653.010 4.280 ;
        RECT 653.850 3.670 656.230 4.280 ;
        RECT 657.070 3.670 659.910 4.280 ;
        RECT 660.750 3.670 663.590 4.280 ;
        RECT 664.430 3.670 666.810 4.280 ;
        RECT 667.650 3.670 670.490 4.280 ;
        RECT 671.330 3.670 674.170 4.280 ;
        RECT 675.010 3.670 677.390 4.280 ;
        RECT 678.230 3.670 681.070 4.280 ;
        RECT 681.910 3.670 684.750 4.280 ;
        RECT 685.590 3.670 687.970 4.280 ;
        RECT 688.810 3.670 691.650 4.280 ;
        RECT 692.490 3.670 695.330 4.280 ;
        RECT 696.170 3.670 698.550 4.280 ;
        RECT 699.390 3.670 702.230 4.280 ;
        RECT 703.070 3.670 705.910 4.280 ;
        RECT 706.750 3.670 709.130 4.280 ;
        RECT 709.970 3.670 712.810 4.280 ;
        RECT 713.650 3.670 716.490 4.280 ;
        RECT 717.330 3.670 719.710 4.280 ;
        RECT 720.550 3.670 723.390 4.280 ;
        RECT 724.230 3.670 727.070 4.280 ;
        RECT 727.910 3.670 730.290 4.280 ;
        RECT 731.130 3.670 733.970 4.280 ;
        RECT 734.810 3.670 737.650 4.280 ;
        RECT 738.490 3.670 740.870 4.280 ;
        RECT 741.710 3.670 744.550 4.280 ;
        RECT 745.390 3.670 748.230 4.280 ;
        RECT 749.070 3.670 751.450 4.280 ;
        RECT 752.290 3.670 755.130 4.280 ;
        RECT 755.970 3.670 758.810 4.280 ;
        RECT 759.650 3.670 762.030 4.280 ;
        RECT 762.870 3.670 765.710 4.280 ;
        RECT 766.550 3.670 769.390 4.280 ;
        RECT 770.230 3.670 772.610 4.280 ;
        RECT 773.450 3.670 776.290 4.280 ;
        RECT 777.130 3.670 779.970 4.280 ;
        RECT 780.810 3.670 783.190 4.280 ;
        RECT 784.030 3.670 786.870 4.280 ;
        RECT 787.710 3.670 790.550 4.280 ;
        RECT 791.390 3.670 793.770 4.280 ;
        RECT 794.610 3.670 797.450 4.280 ;
      LAYER met3 ;
        RECT 4.000 1593.600 795.600 1593.745 ;
        RECT 4.400 1592.880 795.600 1593.600 ;
        RECT 4.400 1592.200 796.000 1592.880 ;
        RECT 4.000 1582.040 796.000 1592.200 ;
        RECT 4.000 1580.640 795.600 1582.040 ;
        RECT 4.000 1580.000 796.000 1580.640 ;
        RECT 4.400 1578.600 796.000 1580.000 ;
        RECT 4.000 1569.800 796.000 1578.600 ;
        RECT 4.000 1568.400 795.600 1569.800 ;
        RECT 4.000 1566.400 796.000 1568.400 ;
        RECT 4.400 1565.000 796.000 1566.400 ;
        RECT 4.000 1557.560 796.000 1565.000 ;
        RECT 4.000 1556.160 795.600 1557.560 ;
        RECT 4.000 1552.800 796.000 1556.160 ;
        RECT 4.400 1551.400 796.000 1552.800 ;
        RECT 4.000 1544.640 796.000 1551.400 ;
        RECT 4.000 1543.240 795.600 1544.640 ;
        RECT 4.000 1539.880 796.000 1543.240 ;
        RECT 4.400 1538.480 796.000 1539.880 ;
        RECT 4.000 1532.400 796.000 1538.480 ;
        RECT 4.000 1531.000 795.600 1532.400 ;
        RECT 4.000 1526.280 796.000 1531.000 ;
        RECT 4.400 1524.880 796.000 1526.280 ;
        RECT 4.000 1520.160 796.000 1524.880 ;
        RECT 4.000 1518.760 795.600 1520.160 ;
        RECT 4.000 1512.680 796.000 1518.760 ;
        RECT 4.400 1511.280 796.000 1512.680 ;
        RECT 4.000 1507.920 796.000 1511.280 ;
        RECT 4.000 1506.520 795.600 1507.920 ;
        RECT 4.000 1499.080 796.000 1506.520 ;
        RECT 4.400 1497.680 796.000 1499.080 ;
        RECT 4.000 1495.000 796.000 1497.680 ;
        RECT 4.000 1493.600 795.600 1495.000 ;
        RECT 4.000 1486.160 796.000 1493.600 ;
        RECT 4.400 1484.760 796.000 1486.160 ;
        RECT 4.000 1482.760 796.000 1484.760 ;
        RECT 4.000 1481.360 795.600 1482.760 ;
        RECT 4.000 1472.560 796.000 1481.360 ;
        RECT 4.400 1471.160 796.000 1472.560 ;
        RECT 4.000 1470.520 796.000 1471.160 ;
        RECT 4.000 1469.120 795.600 1470.520 ;
        RECT 4.000 1458.960 796.000 1469.120 ;
        RECT 4.400 1458.280 796.000 1458.960 ;
        RECT 4.400 1457.560 795.600 1458.280 ;
        RECT 4.000 1456.880 795.600 1457.560 ;
        RECT 4.000 1445.360 796.000 1456.880 ;
        RECT 4.400 1443.960 795.600 1445.360 ;
        RECT 4.000 1433.120 796.000 1443.960 ;
        RECT 4.000 1431.760 795.600 1433.120 ;
        RECT 4.400 1431.720 795.600 1431.760 ;
        RECT 4.400 1430.360 796.000 1431.720 ;
        RECT 4.000 1420.880 796.000 1430.360 ;
        RECT 4.000 1419.480 795.600 1420.880 ;
        RECT 4.000 1418.840 796.000 1419.480 ;
        RECT 4.400 1417.440 796.000 1418.840 ;
        RECT 4.000 1408.640 796.000 1417.440 ;
        RECT 4.000 1407.240 795.600 1408.640 ;
        RECT 4.000 1405.240 796.000 1407.240 ;
        RECT 4.400 1403.840 796.000 1405.240 ;
        RECT 4.000 1395.720 796.000 1403.840 ;
        RECT 4.000 1394.320 795.600 1395.720 ;
        RECT 4.000 1391.640 796.000 1394.320 ;
        RECT 4.400 1390.240 796.000 1391.640 ;
        RECT 4.000 1383.480 796.000 1390.240 ;
        RECT 4.000 1382.080 795.600 1383.480 ;
        RECT 4.000 1378.040 796.000 1382.080 ;
        RECT 4.400 1376.640 796.000 1378.040 ;
        RECT 4.000 1371.240 796.000 1376.640 ;
        RECT 4.000 1369.840 795.600 1371.240 ;
        RECT 4.000 1365.120 796.000 1369.840 ;
        RECT 4.400 1363.720 796.000 1365.120 ;
        RECT 4.000 1359.000 796.000 1363.720 ;
        RECT 4.000 1357.600 795.600 1359.000 ;
        RECT 4.000 1351.520 796.000 1357.600 ;
        RECT 4.400 1350.120 796.000 1351.520 ;
        RECT 4.000 1346.080 796.000 1350.120 ;
        RECT 4.000 1344.680 795.600 1346.080 ;
        RECT 4.000 1337.920 796.000 1344.680 ;
        RECT 4.400 1336.520 796.000 1337.920 ;
        RECT 4.000 1333.840 796.000 1336.520 ;
        RECT 4.000 1332.440 795.600 1333.840 ;
        RECT 4.000 1324.320 796.000 1332.440 ;
        RECT 4.400 1322.920 796.000 1324.320 ;
        RECT 4.000 1321.600 796.000 1322.920 ;
        RECT 4.000 1320.200 795.600 1321.600 ;
        RECT 4.000 1310.720 796.000 1320.200 ;
        RECT 4.400 1309.360 796.000 1310.720 ;
        RECT 4.400 1309.320 795.600 1309.360 ;
        RECT 4.000 1307.960 795.600 1309.320 ;
        RECT 4.000 1297.800 796.000 1307.960 ;
        RECT 4.400 1296.440 796.000 1297.800 ;
        RECT 4.400 1296.400 795.600 1296.440 ;
        RECT 4.000 1295.040 795.600 1296.400 ;
        RECT 4.000 1284.200 796.000 1295.040 ;
        RECT 4.400 1282.800 795.600 1284.200 ;
        RECT 4.000 1271.960 796.000 1282.800 ;
        RECT 4.000 1270.600 795.600 1271.960 ;
        RECT 4.400 1270.560 795.600 1270.600 ;
        RECT 4.400 1269.200 796.000 1270.560 ;
        RECT 4.000 1259.720 796.000 1269.200 ;
        RECT 4.000 1258.320 795.600 1259.720 ;
        RECT 4.000 1257.000 796.000 1258.320 ;
        RECT 4.400 1255.600 796.000 1257.000 ;
        RECT 4.000 1247.480 796.000 1255.600 ;
        RECT 4.000 1246.080 795.600 1247.480 ;
        RECT 4.000 1244.080 796.000 1246.080 ;
        RECT 4.400 1242.680 796.000 1244.080 ;
        RECT 4.000 1234.560 796.000 1242.680 ;
        RECT 4.000 1233.160 795.600 1234.560 ;
        RECT 4.000 1230.480 796.000 1233.160 ;
        RECT 4.400 1229.080 796.000 1230.480 ;
        RECT 4.000 1222.320 796.000 1229.080 ;
        RECT 4.000 1220.920 795.600 1222.320 ;
        RECT 4.000 1216.880 796.000 1220.920 ;
        RECT 4.400 1215.480 796.000 1216.880 ;
        RECT 4.000 1210.080 796.000 1215.480 ;
        RECT 4.000 1208.680 795.600 1210.080 ;
        RECT 4.000 1203.280 796.000 1208.680 ;
        RECT 4.400 1201.880 796.000 1203.280 ;
        RECT 4.000 1197.840 796.000 1201.880 ;
        RECT 4.000 1196.440 795.600 1197.840 ;
        RECT 4.000 1190.360 796.000 1196.440 ;
        RECT 4.400 1188.960 796.000 1190.360 ;
        RECT 4.000 1184.920 796.000 1188.960 ;
        RECT 4.000 1183.520 795.600 1184.920 ;
        RECT 4.000 1176.760 796.000 1183.520 ;
        RECT 4.400 1175.360 796.000 1176.760 ;
        RECT 4.000 1172.680 796.000 1175.360 ;
        RECT 4.000 1171.280 795.600 1172.680 ;
        RECT 4.000 1163.160 796.000 1171.280 ;
        RECT 4.400 1161.760 796.000 1163.160 ;
        RECT 4.000 1160.440 796.000 1161.760 ;
        RECT 4.000 1159.040 795.600 1160.440 ;
        RECT 4.000 1149.560 796.000 1159.040 ;
        RECT 4.400 1148.200 796.000 1149.560 ;
        RECT 4.400 1148.160 795.600 1148.200 ;
        RECT 4.000 1146.800 795.600 1148.160 ;
        RECT 4.000 1135.960 796.000 1146.800 ;
        RECT 4.400 1135.280 796.000 1135.960 ;
        RECT 4.400 1134.560 795.600 1135.280 ;
        RECT 4.000 1133.880 795.600 1134.560 ;
        RECT 4.000 1123.040 796.000 1133.880 ;
        RECT 4.400 1121.640 795.600 1123.040 ;
        RECT 4.000 1110.800 796.000 1121.640 ;
        RECT 4.000 1109.440 795.600 1110.800 ;
        RECT 4.400 1109.400 795.600 1109.440 ;
        RECT 4.400 1108.040 796.000 1109.400 ;
        RECT 4.000 1098.560 796.000 1108.040 ;
        RECT 4.000 1097.160 795.600 1098.560 ;
        RECT 4.000 1095.840 796.000 1097.160 ;
        RECT 4.400 1094.440 796.000 1095.840 ;
        RECT 4.000 1085.640 796.000 1094.440 ;
        RECT 4.000 1084.240 795.600 1085.640 ;
        RECT 4.000 1082.240 796.000 1084.240 ;
        RECT 4.400 1080.840 796.000 1082.240 ;
        RECT 4.000 1073.400 796.000 1080.840 ;
        RECT 4.000 1072.000 795.600 1073.400 ;
        RECT 4.000 1069.320 796.000 1072.000 ;
        RECT 4.400 1067.920 796.000 1069.320 ;
        RECT 4.000 1061.160 796.000 1067.920 ;
        RECT 4.000 1059.760 795.600 1061.160 ;
        RECT 4.000 1055.720 796.000 1059.760 ;
        RECT 4.400 1054.320 796.000 1055.720 ;
        RECT 4.000 1048.920 796.000 1054.320 ;
        RECT 4.000 1047.520 795.600 1048.920 ;
        RECT 4.000 1042.120 796.000 1047.520 ;
        RECT 4.400 1040.720 796.000 1042.120 ;
        RECT 4.000 1036.000 796.000 1040.720 ;
        RECT 4.000 1034.600 795.600 1036.000 ;
        RECT 4.000 1028.520 796.000 1034.600 ;
        RECT 4.400 1027.120 796.000 1028.520 ;
        RECT 4.000 1023.760 796.000 1027.120 ;
        RECT 4.000 1022.360 795.600 1023.760 ;
        RECT 4.000 1014.920 796.000 1022.360 ;
        RECT 4.400 1013.520 796.000 1014.920 ;
        RECT 4.000 1011.520 796.000 1013.520 ;
        RECT 4.000 1010.120 795.600 1011.520 ;
        RECT 4.000 1002.000 796.000 1010.120 ;
        RECT 4.400 1000.600 796.000 1002.000 ;
        RECT 4.000 999.280 796.000 1000.600 ;
        RECT 4.000 997.880 795.600 999.280 ;
        RECT 4.000 988.400 796.000 997.880 ;
        RECT 4.400 987.000 796.000 988.400 ;
        RECT 4.000 986.360 796.000 987.000 ;
        RECT 4.000 984.960 795.600 986.360 ;
        RECT 4.000 974.800 796.000 984.960 ;
        RECT 4.400 974.120 796.000 974.800 ;
        RECT 4.400 973.400 795.600 974.120 ;
        RECT 4.000 972.720 795.600 973.400 ;
        RECT 4.000 961.880 796.000 972.720 ;
        RECT 4.000 961.200 795.600 961.880 ;
        RECT 4.400 960.480 795.600 961.200 ;
        RECT 4.400 959.800 796.000 960.480 ;
        RECT 4.000 949.640 796.000 959.800 ;
        RECT 4.000 948.280 795.600 949.640 ;
        RECT 4.400 948.240 795.600 948.280 ;
        RECT 4.400 946.880 796.000 948.240 ;
        RECT 4.000 937.400 796.000 946.880 ;
        RECT 4.000 936.000 795.600 937.400 ;
        RECT 4.000 934.680 796.000 936.000 ;
        RECT 4.400 933.280 796.000 934.680 ;
        RECT 4.000 924.480 796.000 933.280 ;
        RECT 4.000 923.080 795.600 924.480 ;
        RECT 4.000 921.080 796.000 923.080 ;
        RECT 4.400 919.680 796.000 921.080 ;
        RECT 4.000 912.240 796.000 919.680 ;
        RECT 4.000 910.840 795.600 912.240 ;
        RECT 4.000 907.480 796.000 910.840 ;
        RECT 4.400 906.080 796.000 907.480 ;
        RECT 4.000 900.000 796.000 906.080 ;
        RECT 4.000 898.600 795.600 900.000 ;
        RECT 4.000 894.560 796.000 898.600 ;
        RECT 4.400 893.160 796.000 894.560 ;
        RECT 4.000 887.760 796.000 893.160 ;
        RECT 4.000 886.360 795.600 887.760 ;
        RECT 4.000 880.960 796.000 886.360 ;
        RECT 4.400 879.560 796.000 880.960 ;
        RECT 4.000 874.840 796.000 879.560 ;
        RECT 4.000 873.440 795.600 874.840 ;
        RECT 4.000 867.360 796.000 873.440 ;
        RECT 4.400 865.960 796.000 867.360 ;
        RECT 4.000 862.600 796.000 865.960 ;
        RECT 4.000 861.200 795.600 862.600 ;
        RECT 4.000 853.760 796.000 861.200 ;
        RECT 4.400 852.360 796.000 853.760 ;
        RECT 4.000 850.360 796.000 852.360 ;
        RECT 4.000 848.960 795.600 850.360 ;
        RECT 4.000 840.160 796.000 848.960 ;
        RECT 4.400 838.760 796.000 840.160 ;
        RECT 4.000 838.120 796.000 838.760 ;
        RECT 4.000 836.720 795.600 838.120 ;
        RECT 4.000 827.240 796.000 836.720 ;
        RECT 4.400 825.840 796.000 827.240 ;
        RECT 4.000 825.200 796.000 825.840 ;
        RECT 4.000 823.800 795.600 825.200 ;
        RECT 4.000 813.640 796.000 823.800 ;
        RECT 4.400 812.960 796.000 813.640 ;
        RECT 4.400 812.240 795.600 812.960 ;
        RECT 4.000 811.560 795.600 812.240 ;
        RECT 4.000 800.720 796.000 811.560 ;
        RECT 4.000 800.040 795.600 800.720 ;
        RECT 4.400 799.320 795.600 800.040 ;
        RECT 4.400 798.640 796.000 799.320 ;
        RECT 4.000 788.480 796.000 798.640 ;
        RECT 4.000 787.080 795.600 788.480 ;
        RECT 4.000 786.440 796.000 787.080 ;
        RECT 4.400 785.040 796.000 786.440 ;
        RECT 4.000 775.560 796.000 785.040 ;
        RECT 4.000 774.160 795.600 775.560 ;
        RECT 4.000 773.520 796.000 774.160 ;
        RECT 4.400 772.120 796.000 773.520 ;
        RECT 4.000 763.320 796.000 772.120 ;
        RECT 4.000 761.920 795.600 763.320 ;
        RECT 4.000 759.920 796.000 761.920 ;
        RECT 4.400 758.520 796.000 759.920 ;
        RECT 4.000 751.080 796.000 758.520 ;
        RECT 4.000 749.680 795.600 751.080 ;
        RECT 4.000 746.320 796.000 749.680 ;
        RECT 4.400 744.920 796.000 746.320 ;
        RECT 4.000 738.840 796.000 744.920 ;
        RECT 4.000 737.440 795.600 738.840 ;
        RECT 4.000 732.720 796.000 737.440 ;
        RECT 4.400 731.320 796.000 732.720 ;
        RECT 4.000 725.920 796.000 731.320 ;
        RECT 4.000 724.520 795.600 725.920 ;
        RECT 4.000 719.120 796.000 724.520 ;
        RECT 4.400 717.720 796.000 719.120 ;
        RECT 4.000 713.680 796.000 717.720 ;
        RECT 4.000 712.280 795.600 713.680 ;
        RECT 4.000 706.200 796.000 712.280 ;
        RECT 4.400 704.800 796.000 706.200 ;
        RECT 4.000 701.440 796.000 704.800 ;
        RECT 4.000 700.040 795.600 701.440 ;
        RECT 4.000 692.600 796.000 700.040 ;
        RECT 4.400 691.200 796.000 692.600 ;
        RECT 4.000 689.200 796.000 691.200 ;
        RECT 4.000 687.800 795.600 689.200 ;
        RECT 4.000 679.000 796.000 687.800 ;
        RECT 4.400 677.600 796.000 679.000 ;
        RECT 4.000 676.280 796.000 677.600 ;
        RECT 4.000 674.880 795.600 676.280 ;
        RECT 4.000 665.400 796.000 674.880 ;
        RECT 4.400 664.040 796.000 665.400 ;
        RECT 4.400 664.000 795.600 664.040 ;
        RECT 4.000 662.640 795.600 664.000 ;
        RECT 4.000 652.480 796.000 662.640 ;
        RECT 4.400 651.800 796.000 652.480 ;
        RECT 4.400 651.080 795.600 651.800 ;
        RECT 4.000 650.400 795.600 651.080 ;
        RECT 4.000 639.560 796.000 650.400 ;
        RECT 4.000 638.880 795.600 639.560 ;
        RECT 4.400 638.160 795.600 638.880 ;
        RECT 4.400 637.480 796.000 638.160 ;
        RECT 4.000 627.320 796.000 637.480 ;
        RECT 4.000 625.920 795.600 627.320 ;
        RECT 4.000 625.280 796.000 625.920 ;
        RECT 4.400 623.880 796.000 625.280 ;
        RECT 4.000 614.400 796.000 623.880 ;
        RECT 4.000 613.000 795.600 614.400 ;
        RECT 4.000 611.680 796.000 613.000 ;
        RECT 4.400 610.280 796.000 611.680 ;
        RECT 4.000 602.160 796.000 610.280 ;
        RECT 4.000 600.760 795.600 602.160 ;
        RECT 4.000 598.760 796.000 600.760 ;
        RECT 4.400 597.360 796.000 598.760 ;
        RECT 4.000 589.920 796.000 597.360 ;
        RECT 4.000 588.520 795.600 589.920 ;
        RECT 4.000 585.160 796.000 588.520 ;
        RECT 4.400 583.760 796.000 585.160 ;
        RECT 4.000 577.680 796.000 583.760 ;
        RECT 4.000 576.280 795.600 577.680 ;
        RECT 4.000 571.560 796.000 576.280 ;
        RECT 4.400 570.160 796.000 571.560 ;
        RECT 4.000 564.760 796.000 570.160 ;
        RECT 4.000 563.360 795.600 564.760 ;
        RECT 4.000 557.960 796.000 563.360 ;
        RECT 4.400 556.560 796.000 557.960 ;
        RECT 4.000 552.520 796.000 556.560 ;
        RECT 4.000 551.120 795.600 552.520 ;
        RECT 4.000 544.360 796.000 551.120 ;
        RECT 4.400 542.960 796.000 544.360 ;
        RECT 4.000 540.280 796.000 542.960 ;
        RECT 4.000 538.880 795.600 540.280 ;
        RECT 4.000 531.440 796.000 538.880 ;
        RECT 4.400 530.040 796.000 531.440 ;
        RECT 4.000 528.040 796.000 530.040 ;
        RECT 4.000 526.640 795.600 528.040 ;
        RECT 4.000 517.840 796.000 526.640 ;
        RECT 4.400 516.440 796.000 517.840 ;
        RECT 4.000 515.120 796.000 516.440 ;
        RECT 4.000 513.720 795.600 515.120 ;
        RECT 4.000 504.240 796.000 513.720 ;
        RECT 4.400 502.880 796.000 504.240 ;
        RECT 4.400 502.840 795.600 502.880 ;
        RECT 4.000 501.480 795.600 502.840 ;
        RECT 4.000 490.640 796.000 501.480 ;
        RECT 4.400 489.240 795.600 490.640 ;
        RECT 4.000 478.400 796.000 489.240 ;
        RECT 4.000 477.720 795.600 478.400 ;
        RECT 4.400 477.000 795.600 477.720 ;
        RECT 4.400 476.320 796.000 477.000 ;
        RECT 4.000 465.480 796.000 476.320 ;
        RECT 4.000 464.120 795.600 465.480 ;
        RECT 4.400 464.080 795.600 464.120 ;
        RECT 4.400 462.720 796.000 464.080 ;
        RECT 4.000 453.240 796.000 462.720 ;
        RECT 4.000 451.840 795.600 453.240 ;
        RECT 4.000 450.520 796.000 451.840 ;
        RECT 4.400 449.120 796.000 450.520 ;
        RECT 4.000 441.000 796.000 449.120 ;
        RECT 4.000 439.600 795.600 441.000 ;
        RECT 4.000 436.920 796.000 439.600 ;
        RECT 4.400 435.520 796.000 436.920 ;
        RECT 4.000 428.760 796.000 435.520 ;
        RECT 4.000 427.360 795.600 428.760 ;
        RECT 4.000 423.320 796.000 427.360 ;
        RECT 4.400 421.920 796.000 423.320 ;
        RECT 4.000 415.840 796.000 421.920 ;
        RECT 4.000 414.440 795.600 415.840 ;
        RECT 4.000 410.400 796.000 414.440 ;
        RECT 4.400 409.000 796.000 410.400 ;
        RECT 4.000 403.600 796.000 409.000 ;
        RECT 4.000 402.200 795.600 403.600 ;
        RECT 4.000 396.800 796.000 402.200 ;
        RECT 4.400 395.400 796.000 396.800 ;
        RECT 4.000 391.360 796.000 395.400 ;
        RECT 4.000 389.960 795.600 391.360 ;
        RECT 4.000 383.200 796.000 389.960 ;
        RECT 4.400 381.800 796.000 383.200 ;
        RECT 4.000 379.120 796.000 381.800 ;
        RECT 4.000 377.720 795.600 379.120 ;
        RECT 4.000 369.600 796.000 377.720 ;
        RECT 4.400 368.200 796.000 369.600 ;
        RECT 4.000 366.200 796.000 368.200 ;
        RECT 4.000 364.800 795.600 366.200 ;
        RECT 4.000 356.680 796.000 364.800 ;
        RECT 4.400 355.280 796.000 356.680 ;
        RECT 4.000 353.960 796.000 355.280 ;
        RECT 4.000 352.560 795.600 353.960 ;
        RECT 4.000 343.080 796.000 352.560 ;
        RECT 4.400 341.720 796.000 343.080 ;
        RECT 4.400 341.680 795.600 341.720 ;
        RECT 4.000 340.320 795.600 341.680 ;
        RECT 4.000 329.480 796.000 340.320 ;
        RECT 4.400 328.080 795.600 329.480 ;
        RECT 4.000 317.240 796.000 328.080 ;
        RECT 4.000 315.880 795.600 317.240 ;
        RECT 4.400 315.840 795.600 315.880 ;
        RECT 4.400 314.480 796.000 315.840 ;
        RECT 4.000 304.320 796.000 314.480 ;
        RECT 4.000 302.960 795.600 304.320 ;
        RECT 4.400 302.920 795.600 302.960 ;
        RECT 4.400 301.560 796.000 302.920 ;
        RECT 4.000 292.080 796.000 301.560 ;
        RECT 4.000 290.680 795.600 292.080 ;
        RECT 4.000 289.360 796.000 290.680 ;
        RECT 4.400 287.960 796.000 289.360 ;
        RECT 4.000 279.840 796.000 287.960 ;
        RECT 4.000 278.440 795.600 279.840 ;
        RECT 4.000 275.760 796.000 278.440 ;
        RECT 4.400 274.360 796.000 275.760 ;
        RECT 4.000 267.600 796.000 274.360 ;
        RECT 4.000 266.200 795.600 267.600 ;
        RECT 4.000 262.160 796.000 266.200 ;
        RECT 4.400 260.760 796.000 262.160 ;
        RECT 4.000 254.680 796.000 260.760 ;
        RECT 4.000 253.280 795.600 254.680 ;
        RECT 4.000 248.560 796.000 253.280 ;
        RECT 4.400 247.160 796.000 248.560 ;
        RECT 4.000 242.440 796.000 247.160 ;
        RECT 4.000 241.040 795.600 242.440 ;
        RECT 4.000 235.640 796.000 241.040 ;
        RECT 4.400 234.240 796.000 235.640 ;
        RECT 4.000 230.200 796.000 234.240 ;
        RECT 4.000 228.800 795.600 230.200 ;
        RECT 4.000 222.040 796.000 228.800 ;
        RECT 4.400 220.640 796.000 222.040 ;
        RECT 4.000 217.960 796.000 220.640 ;
        RECT 4.000 216.560 795.600 217.960 ;
        RECT 4.000 208.440 796.000 216.560 ;
        RECT 4.400 207.040 796.000 208.440 ;
        RECT 4.000 205.040 796.000 207.040 ;
        RECT 4.000 203.640 795.600 205.040 ;
        RECT 4.000 194.840 796.000 203.640 ;
        RECT 4.400 193.440 796.000 194.840 ;
        RECT 4.000 192.800 796.000 193.440 ;
        RECT 4.000 191.400 795.600 192.800 ;
        RECT 4.000 181.920 796.000 191.400 ;
        RECT 4.400 180.560 796.000 181.920 ;
        RECT 4.400 180.520 795.600 180.560 ;
        RECT 4.000 179.160 795.600 180.520 ;
        RECT 4.000 168.320 796.000 179.160 ;
        RECT 4.400 166.920 795.600 168.320 ;
        RECT 4.000 155.400 796.000 166.920 ;
        RECT 4.000 154.720 795.600 155.400 ;
        RECT 4.400 154.000 795.600 154.720 ;
        RECT 4.400 153.320 796.000 154.000 ;
        RECT 4.000 143.160 796.000 153.320 ;
        RECT 4.000 141.760 795.600 143.160 ;
        RECT 4.000 141.120 796.000 141.760 ;
        RECT 4.400 139.720 796.000 141.120 ;
        RECT 4.000 130.920 796.000 139.720 ;
        RECT 4.000 129.520 795.600 130.920 ;
        RECT 4.000 127.520 796.000 129.520 ;
        RECT 4.400 126.120 796.000 127.520 ;
        RECT 4.000 118.680 796.000 126.120 ;
        RECT 4.000 117.280 795.600 118.680 ;
        RECT 4.000 114.600 796.000 117.280 ;
        RECT 4.400 113.200 796.000 114.600 ;
        RECT 4.000 105.760 796.000 113.200 ;
        RECT 4.000 104.360 795.600 105.760 ;
        RECT 4.000 101.000 796.000 104.360 ;
        RECT 4.400 99.600 796.000 101.000 ;
        RECT 4.000 93.520 796.000 99.600 ;
        RECT 4.000 92.120 795.600 93.520 ;
        RECT 4.000 87.400 796.000 92.120 ;
        RECT 4.400 86.000 796.000 87.400 ;
        RECT 4.000 81.280 796.000 86.000 ;
        RECT 4.000 79.880 795.600 81.280 ;
        RECT 4.000 73.800 796.000 79.880 ;
        RECT 4.400 72.400 796.000 73.800 ;
        RECT 4.000 69.040 796.000 72.400 ;
        RECT 4.000 67.640 795.600 69.040 ;
        RECT 4.000 60.880 796.000 67.640 ;
        RECT 4.400 59.480 796.000 60.880 ;
        RECT 4.000 56.120 796.000 59.480 ;
        RECT 4.000 54.720 795.600 56.120 ;
        RECT 4.000 47.280 796.000 54.720 ;
        RECT 4.400 45.880 796.000 47.280 ;
        RECT 4.000 43.880 796.000 45.880 ;
        RECT 4.000 42.480 795.600 43.880 ;
        RECT 4.000 33.680 796.000 42.480 ;
        RECT 4.400 32.280 796.000 33.680 ;
        RECT 4.000 31.640 796.000 32.280 ;
        RECT 4.000 30.240 795.600 31.640 ;
        RECT 4.000 20.080 796.000 30.240 ;
        RECT 4.400 19.400 796.000 20.080 ;
        RECT 4.400 18.680 795.600 19.400 ;
        RECT 4.000 18.000 795.600 18.680 ;
        RECT 4.000 7.160 796.000 18.000 ;
        RECT 4.400 6.295 795.600 7.160 ;
      LAYER met4 ;
        RECT 118.055 12.415 174.240 409.185 ;
        RECT 176.640 12.415 239.825 409.185 ;
  END
END user_proj_example
END LIBRARY

