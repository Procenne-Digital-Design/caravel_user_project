module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \sram_addr_a[0] ;
 wire \sram_addr_a[1] ;
 wire \sram_addr_a[2] ;
 wire \sram_addr_a[3] ;
 wire \sram_addr_a[4] ;
 wire \sram_addr_a[5] ;
 wire \sram_addr_a[6] ;
 wire \sram_addr_a[7] ;
 wire \sram_addr_a[8] ;
 wire \sram_addr_b[0] ;
 wire \sram_addr_b[1] ;
 wire \sram_addr_b[2] ;
 wire \sram_addr_b[3] ;
 wire \sram_addr_b[4] ;
 wire \sram_addr_b[5] ;
 wire \sram_addr_b[6] ;
 wire \sram_addr_b[7] ;
 wire \sram_addr_b[8] ;
 wire sram_csb_a;
 wire sram_csb_b;
 wire \sram_din_b[0] ;
 wire \sram_din_b[10] ;
 wire \sram_din_b[11] ;
 wire \sram_din_b[12] ;
 wire \sram_din_b[13] ;
 wire \sram_din_b[14] ;
 wire \sram_din_b[15] ;
 wire \sram_din_b[16] ;
 wire \sram_din_b[17] ;
 wire \sram_din_b[18] ;
 wire \sram_din_b[19] ;
 wire \sram_din_b[1] ;
 wire \sram_din_b[20] ;
 wire \sram_din_b[21] ;
 wire \sram_din_b[22] ;
 wire \sram_din_b[23] ;
 wire \sram_din_b[24] ;
 wire \sram_din_b[25] ;
 wire \sram_din_b[26] ;
 wire \sram_din_b[27] ;
 wire \sram_din_b[28] ;
 wire \sram_din_b[29] ;
 wire \sram_din_b[2] ;
 wire \sram_din_b[30] ;
 wire \sram_din_b[31] ;
 wire \sram_din_b[3] ;
 wire \sram_din_b[4] ;
 wire \sram_din_b[5] ;
 wire \sram_din_b[6] ;
 wire \sram_din_b[7] ;
 wire \sram_din_b[8] ;
 wire \sram_din_b[9] ;
 wire \sram_dout_a[0] ;
 wire \sram_dout_a[10] ;
 wire \sram_dout_a[11] ;
 wire \sram_dout_a[12] ;
 wire \sram_dout_a[13] ;
 wire \sram_dout_a[14] ;
 wire \sram_dout_a[15] ;
 wire \sram_dout_a[16] ;
 wire \sram_dout_a[17] ;
 wire \sram_dout_a[18] ;
 wire \sram_dout_a[19] ;
 wire \sram_dout_a[1] ;
 wire \sram_dout_a[20] ;
 wire \sram_dout_a[21] ;
 wire \sram_dout_a[22] ;
 wire \sram_dout_a[23] ;
 wire \sram_dout_a[24] ;
 wire \sram_dout_a[25] ;
 wire \sram_dout_a[26] ;
 wire \sram_dout_a[27] ;
 wire \sram_dout_a[28] ;
 wire \sram_dout_a[29] ;
 wire \sram_dout_a[2] ;
 wire \sram_dout_a[30] ;
 wire \sram_dout_a[31] ;
 wire \sram_dout_a[3] ;
 wire \sram_dout_a[4] ;
 wire \sram_dout_a[5] ;
 wire \sram_dout_a[6] ;
 wire \sram_dout_a[7] ;
 wire \sram_dout_a[8] ;
 wire \sram_dout_a[9] ;
 wire \sram_mask_b[0] ;
 wire \sram_mask_b[1] ;
 wire \sram_mask_b[2] ;
 wire \sram_mask_b[3] ;
 wire sram_web_b;

 user_proj_example mprj (.sram_csb_a(sram_csb_a),
    .sram_csb_b(sram_csb_b),
    .sram_web_b(sram_web_b),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .io_in({io_in[37],
    io_in[36],
    io_in[35],
    io_in[34],
    io_in[33],
    io_in[32],
    io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21],
    io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .irq({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .la_data_in({la_data_in[127],
    la_data_in[126],
    la_data_in[125],
    la_data_in[124],
    la_data_in[123],
    la_data_in[122],
    la_data_in[121],
    la_data_in[120],
    la_data_in[119],
    la_data_in[118],
    la_data_in[117],
    la_data_in[116],
    la_data_in[115],
    la_data_in[114],
    la_data_in[113],
    la_data_in[112],
    la_data_in[111],
    la_data_in[110],
    la_data_in[109],
    la_data_in[108],
    la_data_in[107],
    la_data_in[106],
    la_data_in[105],
    la_data_in[104],
    la_data_in[103],
    la_data_in[102],
    la_data_in[101],
    la_data_in[100],
    la_data_in[99],
    la_data_in[98],
    la_data_in[97],
    la_data_in[96],
    la_data_in[95],
    la_data_in[94],
    la_data_in[93],
    la_data_in[92],
    la_data_in[91],
    la_data_in[90],
    la_data_in[89],
    la_data_in[88],
    la_data_in[87],
    la_data_in[86],
    la_data_in[85],
    la_data_in[84],
    la_data_in[83],
    la_data_in[82],
    la_data_in[81],
    la_data_in[80],
    la_data_in[79],
    la_data_in[78],
    la_data_in[77],
    la_data_in[76],
    la_data_in[75],
    la_data_in[74],
    la_data_in[73],
    la_data_in[72],
    la_data_in[71],
    la_data_in[70],
    la_data_in[69],
    la_data_in[68],
    la_data_in[67],
    la_data_in[66],
    la_data_in[65],
    la_data_in[64],
    la_data_in[63],
    la_data_in[62],
    la_data_in[61],
    la_data_in[60],
    la_data_in[59],
    la_data_in[58],
    la_data_in[57],
    la_data_in[56],
    la_data_in[55],
    la_data_in[54],
    la_data_in[53],
    la_data_in[52],
    la_data_in[51],
    la_data_in[50],
    la_data_in[49],
    la_data_in[48],
    la_data_in[47],
    la_data_in[46],
    la_data_in[45],
    la_data_in[44],
    la_data_in[43],
    la_data_in[42],
    la_data_in[41],
    la_data_in[40],
    la_data_in[39],
    la_data_in[38],
    la_data_in[37],
    la_data_in[36],
    la_data_in[35],
    la_data_in[34],
    la_data_in[33],
    la_data_in[32],
    la_data_in[31],
    la_data_in[30],
    la_data_in[29],
    la_data_in[28],
    la_data_in[27],
    la_data_in[26],
    la_data_in[25],
    la_data_in[24],
    la_data_in[23],
    la_data_in[22],
    la_data_in[21],
    la_data_in[20],
    la_data_in[19],
    la_data_in[18],
    la_data_in[17],
    la_data_in[16],
    la_data_in[15],
    la_data_in[14],
    la_data_in[13],
    la_data_in[12],
    la_data_in[11],
    la_data_in[10],
    la_data_in[9],
    la_data_in[8],
    la_data_in[7],
    la_data_in[6],
    la_data_in[5],
    la_data_in[4],
    la_data_in[3],
    la_data_in[2],
    la_data_in[1],
    la_data_in[0]}),
    .la_data_out({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96],
    la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64],
    la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .la_oenb({la_oenb[127],
    la_oenb[126],
    la_oenb[125],
    la_oenb[124],
    la_oenb[123],
    la_oenb[122],
    la_oenb[121],
    la_oenb[120],
    la_oenb[119],
    la_oenb[118],
    la_oenb[117],
    la_oenb[116],
    la_oenb[115],
    la_oenb[114],
    la_oenb[113],
    la_oenb[112],
    la_oenb[111],
    la_oenb[110],
    la_oenb[109],
    la_oenb[108],
    la_oenb[107],
    la_oenb[106],
    la_oenb[105],
    la_oenb[104],
    la_oenb[103],
    la_oenb[102],
    la_oenb[101],
    la_oenb[100],
    la_oenb[99],
    la_oenb[98],
    la_oenb[97],
    la_oenb[96],
    la_oenb[95],
    la_oenb[94],
    la_oenb[93],
    la_oenb[92],
    la_oenb[91],
    la_oenb[90],
    la_oenb[89],
    la_oenb[88],
    la_oenb[87],
    la_oenb[86],
    la_oenb[85],
    la_oenb[84],
    la_oenb[83],
    la_oenb[82],
    la_oenb[81],
    la_oenb[80],
    la_oenb[79],
    la_oenb[78],
    la_oenb[77],
    la_oenb[76],
    la_oenb[75],
    la_oenb[74],
    la_oenb[73],
    la_oenb[72],
    la_oenb[71],
    la_oenb[70],
    la_oenb[69],
    la_oenb[68],
    la_oenb[67],
    la_oenb[66],
    la_oenb[65],
    la_oenb[64],
    la_oenb[63],
    la_oenb[62],
    la_oenb[61],
    la_oenb[60],
    la_oenb[59],
    la_oenb[58],
    la_oenb[57],
    la_oenb[56],
    la_oenb[55],
    la_oenb[54],
    la_oenb[53],
    la_oenb[52],
    la_oenb[51],
    la_oenb[50],
    la_oenb[49],
    la_oenb[48],
    la_oenb[47],
    la_oenb[46],
    la_oenb[45],
    la_oenb[44],
    la_oenb[43],
    la_oenb[42],
    la_oenb[41],
    la_oenb[40],
    la_oenb[39],
    la_oenb[38],
    la_oenb[37],
    la_oenb[36],
    la_oenb[35],
    la_oenb[34],
    la_oenb[33],
    la_oenb[32],
    la_oenb[31],
    la_oenb[30],
    la_oenb[29],
    la_oenb[28],
    la_oenb[27],
    la_oenb[26],
    la_oenb[25],
    la_oenb[24],
    la_oenb[23],
    la_oenb[22],
    la_oenb[21],
    la_oenb[20],
    la_oenb[19],
    la_oenb[18],
    la_oenb[17],
    la_oenb[16],
    la_oenb[15],
    la_oenb[14],
    la_oenb[13],
    la_oenb[12],
    la_oenb[11],
    la_oenb[10],
    la_oenb[9],
    la_oenb[8],
    la_oenb[7],
    la_oenb[6],
    la_oenb[5],
    la_oenb[4],
    la_oenb[3],
    la_oenb[2],
    la_oenb[1],
    la_oenb[0]}),
    .sram_addr_a({\sram_addr_a[8] ,
    \sram_addr_a[7] ,
    \sram_addr_a[6] ,
    \sram_addr_a[5] ,
    \sram_addr_a[4] ,
    \sram_addr_a[3] ,
    \sram_addr_a[2] ,
    \sram_addr_a[1] ,
    \sram_addr_a[0] }),
    .sram_addr_b({\sram_addr_b[8] ,
    \sram_addr_b[7] ,
    \sram_addr_b[6] ,
    \sram_addr_b[5] ,
    \sram_addr_b[4] ,
    \sram_addr_b[3] ,
    \sram_addr_b[2] ,
    \sram_addr_b[1] ,
    \sram_addr_b[0] }),
    .sram_din_b({\sram_din_b[31] ,
    \sram_din_b[30] ,
    \sram_din_b[29] ,
    \sram_din_b[28] ,
    \sram_din_b[27] ,
    \sram_din_b[26] ,
    \sram_din_b[25] ,
    \sram_din_b[24] ,
    \sram_din_b[23] ,
    \sram_din_b[22] ,
    \sram_din_b[21] ,
    \sram_din_b[20] ,
    \sram_din_b[19] ,
    \sram_din_b[18] ,
    \sram_din_b[17] ,
    \sram_din_b[16] ,
    \sram_din_b[15] ,
    \sram_din_b[14] ,
    \sram_din_b[13] ,
    \sram_din_b[12] ,
    \sram_din_b[11] ,
    \sram_din_b[10] ,
    \sram_din_b[9] ,
    \sram_din_b[8] ,
    \sram_din_b[7] ,
    \sram_din_b[6] ,
    \sram_din_b[5] ,
    \sram_din_b[4] ,
    \sram_din_b[3] ,
    \sram_din_b[2] ,
    \sram_din_b[1] ,
    \sram_din_b[0] }),
    .sram_dout_a({\sram_dout_a[31] ,
    \sram_dout_a[30] ,
    \sram_dout_a[29] ,
    \sram_dout_a[28] ,
    \sram_dout_a[27] ,
    \sram_dout_a[26] ,
    \sram_dout_a[25] ,
    \sram_dout_a[24] ,
    \sram_dout_a[23] ,
    \sram_dout_a[22] ,
    \sram_dout_a[21] ,
    \sram_dout_a[20] ,
    \sram_dout_a[19] ,
    \sram_dout_a[18] ,
    \sram_dout_a[17] ,
    \sram_dout_a[16] ,
    \sram_dout_a[15] ,
    \sram_dout_a[14] ,
    \sram_dout_a[13] ,
    \sram_dout_a[12] ,
    \sram_dout_a[11] ,
    \sram_dout_a[10] ,
    \sram_dout_a[9] ,
    \sram_dout_a[8] ,
    \sram_dout_a[7] ,
    \sram_dout_a[6] ,
    \sram_dout_a[5] ,
    \sram_dout_a[4] ,
    \sram_dout_a[3] ,
    \sram_dout_a[2] ,
    \sram_dout_a[1] ,
    \sram_dout_a[0] }),
    .sram_mask_b({\sram_mask_b[3] ,
    \sram_mask_b[2] ,
    \sram_mask_b[1] ,
    \sram_mask_b[0] }),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 sky130_sram_2kbyte_1rw1r_32x512_8 u_sram1_2kb (.csb0(sram_csb_b),
    .csb1(sram_csb_a),
    .web0(sram_web_b),
    .clk0(wb_clk_i),
    .clk1(wb_clk_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\sram_addr_b[8] ,
    \sram_addr_b[7] ,
    \sram_addr_b[6] ,
    \sram_addr_b[5] ,
    \sram_addr_b[4] ,
    \sram_addr_b[3] ,
    \sram_addr_b[2] ,
    \sram_addr_b[1] ,
    \sram_addr_b[0] }),
    .addr1({\sram_addr_a[8] ,
    \sram_addr_a[7] ,
    \sram_addr_a[6] ,
    \sram_addr_a[5] ,
    \sram_addr_a[4] ,
    \sram_addr_a[3] ,
    \sram_addr_a[2] ,
    \sram_addr_a[1] ,
    \sram_addr_a[0] }),
    .din0({\sram_din_b[31] ,
    \sram_din_b[30] ,
    \sram_din_b[29] ,
    \sram_din_b[28] ,
    \sram_din_b[27] ,
    \sram_din_b[26] ,
    \sram_din_b[25] ,
    \sram_din_b[24] ,
    \sram_din_b[23] ,
    \sram_din_b[22] ,
    \sram_din_b[21] ,
    \sram_din_b[20] ,
    \sram_din_b[19] ,
    \sram_din_b[18] ,
    \sram_din_b[17] ,
    \sram_din_b[16] ,
    \sram_din_b[15] ,
    \sram_din_b[14] ,
    \sram_din_b[13] ,
    \sram_din_b[12] ,
    \sram_din_b[11] ,
    \sram_din_b[10] ,
    \sram_din_b[9] ,
    \sram_din_b[8] ,
    \sram_din_b[7] ,
    \sram_din_b[6] ,
    \sram_din_b[5] ,
    \sram_din_b[4] ,
    \sram_din_b[3] ,
    \sram_din_b[2] ,
    \sram_din_b[1] ,
    \sram_din_b[0] }),
    .dout0({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .dout1({\sram_dout_a[31] ,
    \sram_dout_a[30] ,
    \sram_dout_a[29] ,
    \sram_dout_a[28] ,
    \sram_dout_a[27] ,
    \sram_dout_a[26] ,
    \sram_dout_a[25] ,
    \sram_dout_a[24] ,
    \sram_dout_a[23] ,
    \sram_dout_a[22] ,
    \sram_dout_a[21] ,
    \sram_dout_a[20] ,
    \sram_dout_a[19] ,
    \sram_dout_a[18] ,
    \sram_dout_a[17] ,
    \sram_dout_a[16] ,
    \sram_dout_a[15] ,
    \sram_dout_a[14] ,
    \sram_dout_a[13] ,
    \sram_dout_a[12] ,
    \sram_dout_a[11] ,
    \sram_dout_a[10] ,
    \sram_dout_a[9] ,
    \sram_dout_a[8] ,
    \sram_dout_a[7] ,
    \sram_dout_a[6] ,
    \sram_dout_a[5] ,
    \sram_dout_a[4] ,
    \sram_dout_a[3] ,
    \sram_dout_a[2] ,
    \sram_dout_a[1] ,
    \sram_dout_a[0] }),
    .wmask0({\sram_mask_b[3] ,
    \sram_mask_b[2] ,
    \sram_mask_b[1] ,
    \sram_mask_b[0] }));
endmodule
