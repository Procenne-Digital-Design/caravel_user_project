VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 1600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 1596.000 1.750 1600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1596.000 103.410 1600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 1596.000 113.530 1600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 1596.000 123.650 1600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 1596.000 133.770 1600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 1596.000 143.890 1600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 1596.000 154.010 1600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 1596.000 164.130 1600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1596.000 174.250 1600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 1596.000 184.370 1600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 1596.000 194.950 1600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 1596.000 11.870 1600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 1596.000 205.070 1600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 1596.000 215.190 1600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 1596.000 225.310 1600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1596.000 235.430 1600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 1596.000 245.550 1600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 1596.000 255.670 1600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 1596.000 265.790 1600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 1596.000 275.910 1600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 1596.000 286.030 1600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 1596.000 296.610 1600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 1596.000 21.990 1600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 1596.000 306.730 1600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 1596.000 316.850 1600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 1596.000 326.970 1600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 1596.000 337.090 1600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 1596.000 347.210 1600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 1596.000 357.330 1600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1596.000 367.450 1600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 1596.000 377.570 1600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 1596.000 32.110 1600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1596.000 42.230 1600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 1596.000 52.350 1600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 1596.000 62.470 1600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 1596.000 72.590 1600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 1596.000 82.710 1600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 1596.000 92.830 1600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 1596.000 4.970 1600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 1596.000 106.630 1600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 1596.000 116.750 1600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 1596.000 126.870 1600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 1596.000 136.990 1600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 1596.000 147.110 1600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 1596.000 157.230 1600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1596.000 167.810 1600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 1596.000 177.930 1600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 1596.000 188.050 1600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 1596.000 198.170 1600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 1596.000 15.090 1600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 1596.000 208.290 1600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 1596.000 218.410 1600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 1596.000 228.530 1600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 1596.000 238.650 1600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 1596.000 248.770 1600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 1596.000 259.350 1600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 1596.000 269.470 1600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 1596.000 279.590 1600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 1596.000 289.710 1600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1596.000 299.830 1600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 1596.000 25.210 1600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 1596.000 309.950 1600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 1596.000 320.070 1600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 1596.000 330.190 1600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 1596.000 340.310 1600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 1596.000 350.430 1600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 1596.000 361.010 1600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 1596.000 371.130 1600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 1596.000 381.250 1600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 1596.000 35.330 1600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1596.000 45.450 1600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 1596.000 55.570 1600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 1596.000 66.150 1600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 1596.000 76.270 1600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 1596.000 86.390 1600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 1596.000 96.510 1600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1596.000 8.190 1600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1596.000 109.850 1600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 1596.000 119.970 1600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 1596.000 130.550 1600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 1596.000 140.670 1600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 1596.000 150.790 1600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 1596.000 160.910 1600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1596.000 171.030 1600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 1596.000 181.150 1600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 1596.000 191.270 1600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 1596.000 201.390 1600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 1596.000 18.310 1600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 1596.000 211.510 1600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 1596.000 221.630 1600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 1596.000 232.210 1600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 1596.000 242.330 1600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 1596.000 252.450 1600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 1596.000 262.570 1600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 1596.000 272.690 1600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 1596.000 282.810 1600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 1596.000 292.930 1600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 1596.000 303.050 1600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 1596.000 28.430 1600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 1596.000 313.170 1600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 1596.000 323.750 1600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 1596.000 333.870 1600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 1596.000 343.990 1600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 1596.000 354.110 1600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1596.000 364.230 1600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 1596.000 374.350 1600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 1596.000 384.470 1600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1596.000 39.010 1600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 1596.000 49.130 1600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 1596.000 59.250 1600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 1596.000 69.370 1600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 1596.000 79.490 1600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 1596.000 89.610 1600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 1596.000 99.730 1600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 1596.000 720.270 1600.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.200 4.000 1300.800 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 1596.000 736.830 1600.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1457.280 800.000 1457.880 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 0.000 757.990 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 1596.000 462.670 1600.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1596.000 747.410 1600.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.960 4.000 1356.560 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1487.200 800.000 1487.800 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1502.160 800.000 1502.760 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.120 4.000 1398.720 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1426.000 4.000 1426.600 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1439.600 4.000 1440.200 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 1596.000 763.970 1600.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1453.200 4.000 1453.800 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 395.120 800.000 395.720 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 1596.000 777.770 1600.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1495.360 4.000 1495.960 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 1596.000 784.670 1600.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 1596.000 791.110 1600.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1551.120 4.000 1551.720 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1592.600 4.000 1593.200 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 425.040 800.000 425.640 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 1596.000 479.230 1600.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 1596.000 496.250 1600.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 1596.000 503.150 1600.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 80.960 800.000 81.560 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 1596.000 513.270 1600.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 559.680 800.000 560.280 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 574.640 800.000 575.240 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 1596.000 537.190 1600.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 1596.000 543.630 1600.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 110.880 800.000 111.480 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 604.560 800.000 605.160 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 634.480 800.000 635.080 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 664.400 800.000 665.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 1596.000 574.450 1600.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 1596.000 584.570 1600.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 799.040 800.000 799.640 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 1596.000 591.470 1600.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 828.960 800.000 829.560 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 858.880 800.000 859.480 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 1596.000 597.910 1600.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 1596.000 601.590 1600.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 1596.000 611.710 1600.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 230.560 800.000 231.160 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.720 4.000 953.320 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 966.320 4.000 966.920 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 948.640 800.000 949.240 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1596.000 625.050 1600.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 1596.000 628.730 1600.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 305.360 800.000 305.960 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 993.520 800.000 994.120 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 1596.000 638.850 1600.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 1596.000 642.070 1600.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 1596.000 645.750 1600.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 1596.000 652.190 1600.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1038.400 800.000 1039.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1068.320 800.000 1068.920 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1098.240 800.000 1098.840 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1113.200 800.000 1113.800 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.720 4.000 1106.320 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 1596.000 672.430 1600.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1173.040 800.000 1173.640 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1119.320 4.000 1119.920 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 1596.000 686.230 1600.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1202.960 800.000 1203.560 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 1596.000 445.650 1600.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1232.880 800.000 1233.480 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1247.840 800.000 1248.440 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1277.760 800.000 1278.360 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1189.360 4.000 1189.960 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1322.640 800.000 1323.240 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1367.520 800.000 1368.120 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1382.480 800.000 1383.080 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1272.320 4.000 1272.920 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 1596.000 452.550 1600.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 1596.000 388.150 1600.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1412.400 800.000 1413.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 1596.000 716.590 1600.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 1596.000 723.490 1600.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1286.600 4.000 1287.200 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 1596.000 740.510 1600.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1442.320 800.000 1442.920 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1328.080 4.000 1328.680 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 0.000 761.210 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 365.200 800.000 365.800 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1596.000 753.850 1600.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1517.120 800.000 1517.720 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1532.080 800.000 1532.680 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 1596.000 757.530 1600.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 1596.000 767.650 1600.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1467.480 4.000 1468.080 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 1596.000 469.110 1600.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1481.080 4.000 1481.680 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 1596.000 780.990 1600.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 1596.000 787.890 1600.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1576.960 800.000 1577.560 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 1596.000 794.790 1600.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1579.000 4.000 1579.600 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 1596.000 476.010 1600.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 1596.000 486.130 1600.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 544.720 800.000 545.320 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 1596.000 520.170 1600.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 1596.000 527.070 1600.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 1596.000 540.410 1600.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 1596.000 398.270 1600.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 649.440 800.000 650.040 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1596.000 560.650 1600.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 679.360 800.000 679.960 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 1596.000 570.770 1600.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 170.720 800.000 171.320 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 709.280 800.000 709.880 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 1596.000 577.670 1600.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 1596.000 581.350 1600.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 754.160 800.000 754.760 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 769.120 800.000 769.720 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 1596.000 408.390 1600.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 1596.000 587.790 1600.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.200 4.000 841.800 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 1596.000 594.690 1600.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 873.840 800.000 874.440 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 1596.000 608.030 1600.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 245.520 800.000 246.120 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 903.760 800.000 904.360 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 963.600 800.000 964.200 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1008.480 4.000 1009.080 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 978.560 800.000 979.160 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.960 4.000 1050.560 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1008.480 800.000 1009.080 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 1596.000 655.870 1600.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1083.280 800.000 1083.880 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 335.280 800.000 335.880 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 1596.000 665.990 1600.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1128.160 800.000 1128.760 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1143.120 800.000 1143.720 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 1596.000 676.110 1600.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 1596.000 679.330 1600.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1188.000 800.000 1188.600 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1596.000 689.450 1600.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.200 4.000 1147.800 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 1596.000 693.130 1600.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1262.800 800.000 1263.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 1596.000 699.570 1600.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.960 4.000 1203.560 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1337.600 800.000 1338.200 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 1596.000 703.250 1600.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.120 4.000 1245.720 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 1596.000 710.150 1600.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1397.440 800.000 1398.040 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 1596.000 455.770 1600.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 1596.000 713.370 1600.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 1596.000 726.710 1600.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 1596.000 730.390 1600.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 1596.000 733.610 1600.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1427.360 800.000 1427.960 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 1596.000 743.730 1600.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 4.000 1342.960 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 380.160 800.000 380.760 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1472.240 800.000 1472.840 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 1596.000 750.630 1600.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.720 4.000 1412.320 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1547.040 800.000 1547.640 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 1596.000 760.750 1600.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 1596.000 770.870 1600.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 0.000 774.550 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 1596.000 774.550 1600.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 1596.000 472.790 1600.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1562.000 800.000 1562.600 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1508.960 4.000 1509.560 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 0.000 784.670 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1591.920 800.000 1592.520 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.720 4.000 1565.320 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 1596.000 798.010 1600.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1596.000 489.810 1600.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 1596.000 394.590 1600.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 1596.000 510.050 1600.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 514.800 800.000 515.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 1596.000 523.390 1600.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 589.600 800.000 590.200 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 125.840 800.000 126.440 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 1596.000 547.310 1600.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 619.520 800.000 620.120 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 1596.000 554.210 1600.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 1596.000 557.430 1600.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 1596.000 564.330 1600.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 1596.000 567.550 1600.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 694.320 800.000 694.920 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 1596.000 401.490 1600.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 724.240 800.000 724.840 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 739.200 800.000 739.800 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 784.080 800.000 784.680 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 827.600 4.000 828.200 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 1596.000 411.610 1600.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 814.000 800.000 814.600 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 843.920 800.000 844.520 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.080 4.000 869.680 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 883.360 4.000 883.960 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1596.000 604.810 1600.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 888.800 800.000 889.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 260.480 800.000 261.080 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 910.560 4.000 911.160 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 1596.000 614.930 1600.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 1596.000 618.610 1600.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 918.720 800.000 919.320 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 933.680 800.000 934.280 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1596.000 621.830 1600.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 1596.000 631.950 1600.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 1596.000 425.410 1600.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.080 4.000 1022.680 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 1596.000 635.170 1600.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 1596.000 648.970 1600.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1023.440 800.000 1024.040 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1053.360 800.000 1053.960 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 1596.000 659.090 1600.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 1596.000 662.310 1600.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 1596.000 435.530 1600.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 1596.000 669.210 1600.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1158.080 800.000 1158.680 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1596.000 683.010 1600.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1133.600 4.000 1134.200 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1217.920 800.000 1218.520 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 1596.000 696.350 1600.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1161.480 4.000 1162.080 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1175.080 4.000 1175.680 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1292.720 800.000 1293.320 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1307.680 800.000 1308.280 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1352.560 800.000 1353.160 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 1596.000 706.470 1600.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.720 4.000 1259.320 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END la_oenb[9]
  PIN sram_addr_a[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 36.080 800.000 36.680 ;
    END
  END sram_addr_a[0]
  PIN sram_addr_a[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END sram_addr_a[1]
  PIN sram_addr_a[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END sram_addr_a[2]
  PIN sram_addr_a[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END sram_addr_a[3]
  PIN sram_addr_a[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 200.640 800.000 201.240 ;
    END
  END sram_addr_a[4]
  PIN sram_addr_a[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 275.440 800.000 276.040 ;
    END
  END sram_addr_a[5]
  PIN sram_addr_a[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1596.000 428.630 1600.000 ;
    END
  END sram_addr_a[6]
  PIN sram_addr_a[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 1596.000 438.750 1600.000 ;
    END
  END sram_addr_a[7]
  PIN sram_addr_a[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 1596.000 448.870 1600.000 ;
    END
  END sram_addr_a[8]
  PIN sram_addr_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 51.040 800.000 51.640 ;
    END
  END sram_addr_b[0]
  PIN sram_addr_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END sram_addr_b[1]
  PIN sram_addr_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 140.800 800.000 141.400 ;
    END
  END sram_addr_b[2]
  PIN sram_addr_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 185.680 800.000 186.280 ;
    END
  END sram_addr_b[3]
  PIN sram_addr_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 1596.000 414.830 1600.000 ;
    END
  END sram_addr_b[4]
  PIN sram_addr_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END sram_addr_b[5]
  PIN sram_addr_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 320.320 800.000 320.920 ;
    END
  END sram_addr_b[6]
  PIN sram_addr_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END sram_addr_b[7]
  PIN sram_addr_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 350.240 800.000 350.840 ;
    END
  END sram_addr_b[8]
  PIN sram_csb_a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 6.840 800.000 7.440 ;
    END
  END sram_csb_a
  PIN sram_csb_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END sram_csb_b
  PIN sram_din_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END sram_din_b[0]
  PIN sram_din_b[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END sram_din_b[10]
  PIN sram_din_b[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 410.080 800.000 410.680 ;
    END
  END sram_din_b[11]
  PIN sram_din_b[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 440.000 800.000 440.600 ;
    END
  END sram_din_b[12]
  PIN sram_din_b[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END sram_din_b[13]
  PIN sram_din_b[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END sram_din_b[14]
  PIN sram_din_b[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END sram_din_b[15]
  PIN sram_din_b[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END sram_din_b[16]
  PIN sram_din_b[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 1596.000 499.930 1600.000 ;
    END
  END sram_din_b[17]
  PIN sram_din_b[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END sram_din_b[18]
  PIN sram_din_b[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END sram_din_b[19]
  PIN sram_din_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END sram_din_b[1]
  PIN sram_din_b[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 484.880 800.000 485.480 ;
    END
  END sram_din_b[20]
  PIN sram_din_b[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 529.760 800.000 530.360 ;
    END
  END sram_din_b[21]
  PIN sram_din_b[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END sram_din_b[22]
  PIN sram_din_b[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END sram_din_b[23]
  PIN sram_din_b[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 1596.000 530.290 1600.000 ;
    END
  END sram_din_b[24]
  PIN sram_din_b[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END sram_din_b[25]
  PIN sram_din_b[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 1596.000 533.510 1600.000 ;
    END
  END sram_din_b[26]
  PIN sram_din_b[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END sram_din_b[27]
  PIN sram_din_b[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END sram_din_b[28]
  PIN sram_din_b[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END sram_din_b[29]
  PIN sram_din_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END sram_din_b[2]
  PIN sram_din_b[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END sram_din_b[30]
  PIN sram_din_b[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END sram_din_b[31]
  PIN sram_din_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END sram_din_b[3]
  PIN sram_din_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 1596.000 418.510 1600.000 ;
    END
  END sram_din_b[4]
  PIN sram_din_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 1596.000 421.730 1600.000 ;
    END
  END sram_din_b[5]
  PIN sram_din_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 1596.000 431.850 1600.000 ;
    END
  END sram_din_b[6]
  PIN sram_din_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 1596.000 441.970 1600.000 ;
    END
  END sram_din_b[7]
  PIN sram_din_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END sram_din_b[8]
  PIN sram_din_b[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END sram_din_b[9]
  PIN sram_dout_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 1596.000 391.370 1600.000 ;
    END
  END sram_dout_a[0]
  PIN sram_dout_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 1596.000 465.890 1600.000 ;
    END
  END sram_dout_a[10]
  PIN sram_dout_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END sram_dout_a[11]
  PIN sram_dout_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END sram_dout_a[12]
  PIN sram_dout_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END sram_dout_a[13]
  PIN sram_dout_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 1596.000 482.910 1600.000 ;
    END
  END sram_dout_a[14]
  PIN sram_dout_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 454.960 800.000 455.560 ;
    END
  END sram_dout_a[15]
  PIN sram_dout_a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 1596.000 493.030 1600.000 ;
    END
  END sram_dout_a[16]
  PIN sram_dout_a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END sram_dout_a[17]
  PIN sram_dout_a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 469.920 800.000 470.520 ;
    END
  END sram_dout_a[18]
  PIN sram_dout_a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 1596.000 506.370 1600.000 ;
    END
  END sram_dout_a[19]
  PIN sram_dout_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END sram_dout_a[1]
  PIN sram_dout_a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 499.840 800.000 500.440 ;
    END
  END sram_dout_a[20]
  PIN sram_dout_a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END sram_dout_a[21]
  PIN sram_dout_a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 1596.000 516.950 1600.000 ;
    END
  END sram_dout_a[22]
  PIN sram_dout_a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END sram_dout_a[23]
  PIN sram_dout_a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END sram_dout_a[24]
  PIN sram_dout_a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END sram_dout_a[25]
  PIN sram_dout_a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END sram_dout_a[26]
  PIN sram_dout_a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END sram_dout_a[27]
  PIN sram_dout_a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 521.600 4.000 522.200 ;
    END
  END sram_dout_a[28]
  PIN sram_dout_a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END sram_dout_a[29]
  PIN sram_dout_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END sram_dout_a[2]
  PIN sram_dout_a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END sram_dout_a[30]
  PIN sram_dout_a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 1596.000 550.530 1600.000 ;
    END
  END sram_dout_a[31]
  PIN sram_dout_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END sram_dout_a[3]
  PIN sram_dout_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 215.600 800.000 216.200 ;
    END
  END sram_dout_a[4]
  PIN sram_dout_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 290.400 800.000 291.000 ;
    END
  END sram_dout_a[5]
  PIN sram_dout_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END sram_dout_a[6]
  PIN sram_dout_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END sram_dout_a[7]
  PIN sram_dout_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END sram_dout_a[8]
  PIN sram_dout_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 1596.000 458.990 1600.000 ;
    END
  END sram_dout_a[9]
  PIN sram_mask_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 66.000 800.000 66.600 ;
    END
  END sram_mask_b[0]
  PIN sram_mask_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 95.920 800.000 96.520 ;
    END
  END sram_mask_b[1]
  PIN sram_mask_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 155.760 800.000 156.360 ;
    END
  END sram_mask_b[2]
  PIN sram_mask_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 1596.000 404.710 1600.000 ;
    END
  END sram_mask_b[3]
  PIN sram_web_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 21.120 800.000 21.720 ;
    END
  END sram_web_b
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1588.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1588.720 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 1588.565 ;
      LAYER met1 ;
        RECT 0.070 5.480 794.810 1591.500 ;
      LAYER met2 ;
        RECT 0.100 1595.720 1.190 1596.370 ;
        RECT 2.030 1595.720 4.410 1596.370 ;
        RECT 5.250 1595.720 7.630 1596.370 ;
        RECT 8.470 1595.720 11.310 1596.370 ;
        RECT 12.150 1595.720 14.530 1596.370 ;
        RECT 15.370 1595.720 17.750 1596.370 ;
        RECT 18.590 1595.720 21.430 1596.370 ;
        RECT 22.270 1595.720 24.650 1596.370 ;
        RECT 25.490 1595.720 27.870 1596.370 ;
        RECT 28.710 1595.720 31.550 1596.370 ;
        RECT 32.390 1595.720 34.770 1596.370 ;
        RECT 35.610 1595.720 38.450 1596.370 ;
        RECT 39.290 1595.720 41.670 1596.370 ;
        RECT 42.510 1595.720 44.890 1596.370 ;
        RECT 45.730 1595.720 48.570 1596.370 ;
        RECT 49.410 1595.720 51.790 1596.370 ;
        RECT 52.630 1595.720 55.010 1596.370 ;
        RECT 55.850 1595.720 58.690 1596.370 ;
        RECT 59.530 1595.720 61.910 1596.370 ;
        RECT 62.750 1595.720 65.590 1596.370 ;
        RECT 66.430 1595.720 68.810 1596.370 ;
        RECT 69.650 1595.720 72.030 1596.370 ;
        RECT 72.870 1595.720 75.710 1596.370 ;
        RECT 76.550 1595.720 78.930 1596.370 ;
        RECT 79.770 1595.720 82.150 1596.370 ;
        RECT 82.990 1595.720 85.830 1596.370 ;
        RECT 86.670 1595.720 89.050 1596.370 ;
        RECT 89.890 1595.720 92.270 1596.370 ;
        RECT 93.110 1595.720 95.950 1596.370 ;
        RECT 96.790 1595.720 99.170 1596.370 ;
        RECT 100.010 1595.720 102.850 1596.370 ;
        RECT 103.690 1595.720 106.070 1596.370 ;
        RECT 106.910 1595.720 109.290 1596.370 ;
        RECT 110.130 1595.720 112.970 1596.370 ;
        RECT 113.810 1595.720 116.190 1596.370 ;
        RECT 117.030 1595.720 119.410 1596.370 ;
        RECT 120.250 1595.720 123.090 1596.370 ;
        RECT 123.930 1595.720 126.310 1596.370 ;
        RECT 127.150 1595.720 129.990 1596.370 ;
        RECT 130.830 1595.720 133.210 1596.370 ;
        RECT 134.050 1595.720 136.430 1596.370 ;
        RECT 137.270 1595.720 140.110 1596.370 ;
        RECT 140.950 1595.720 143.330 1596.370 ;
        RECT 144.170 1595.720 146.550 1596.370 ;
        RECT 147.390 1595.720 150.230 1596.370 ;
        RECT 151.070 1595.720 153.450 1596.370 ;
        RECT 154.290 1595.720 156.670 1596.370 ;
        RECT 157.510 1595.720 160.350 1596.370 ;
        RECT 161.190 1595.720 163.570 1596.370 ;
        RECT 164.410 1595.720 167.250 1596.370 ;
        RECT 168.090 1595.720 170.470 1596.370 ;
        RECT 171.310 1595.720 173.690 1596.370 ;
        RECT 174.530 1595.720 177.370 1596.370 ;
        RECT 178.210 1595.720 180.590 1596.370 ;
        RECT 181.430 1595.720 183.810 1596.370 ;
        RECT 184.650 1595.720 187.490 1596.370 ;
        RECT 188.330 1595.720 190.710 1596.370 ;
        RECT 191.550 1595.720 194.390 1596.370 ;
        RECT 195.230 1595.720 197.610 1596.370 ;
        RECT 198.450 1595.720 200.830 1596.370 ;
        RECT 201.670 1595.720 204.510 1596.370 ;
        RECT 205.350 1595.720 207.730 1596.370 ;
        RECT 208.570 1595.720 210.950 1596.370 ;
        RECT 211.790 1595.720 214.630 1596.370 ;
        RECT 215.470 1595.720 217.850 1596.370 ;
        RECT 218.690 1595.720 221.070 1596.370 ;
        RECT 221.910 1595.720 224.750 1596.370 ;
        RECT 225.590 1595.720 227.970 1596.370 ;
        RECT 228.810 1595.720 231.650 1596.370 ;
        RECT 232.490 1595.720 234.870 1596.370 ;
        RECT 235.710 1595.720 238.090 1596.370 ;
        RECT 238.930 1595.720 241.770 1596.370 ;
        RECT 242.610 1595.720 244.990 1596.370 ;
        RECT 245.830 1595.720 248.210 1596.370 ;
        RECT 249.050 1595.720 251.890 1596.370 ;
        RECT 252.730 1595.720 255.110 1596.370 ;
        RECT 255.950 1595.720 258.790 1596.370 ;
        RECT 259.630 1595.720 262.010 1596.370 ;
        RECT 262.850 1595.720 265.230 1596.370 ;
        RECT 266.070 1595.720 268.910 1596.370 ;
        RECT 269.750 1595.720 272.130 1596.370 ;
        RECT 272.970 1595.720 275.350 1596.370 ;
        RECT 276.190 1595.720 279.030 1596.370 ;
        RECT 279.870 1595.720 282.250 1596.370 ;
        RECT 283.090 1595.720 285.470 1596.370 ;
        RECT 286.310 1595.720 289.150 1596.370 ;
        RECT 289.990 1595.720 292.370 1596.370 ;
        RECT 293.210 1595.720 296.050 1596.370 ;
        RECT 296.890 1595.720 299.270 1596.370 ;
        RECT 300.110 1595.720 302.490 1596.370 ;
        RECT 303.330 1595.720 306.170 1596.370 ;
        RECT 307.010 1595.720 309.390 1596.370 ;
        RECT 310.230 1595.720 312.610 1596.370 ;
        RECT 313.450 1595.720 316.290 1596.370 ;
        RECT 317.130 1595.720 319.510 1596.370 ;
        RECT 320.350 1595.720 323.190 1596.370 ;
        RECT 324.030 1595.720 326.410 1596.370 ;
        RECT 327.250 1595.720 329.630 1596.370 ;
        RECT 330.470 1595.720 333.310 1596.370 ;
        RECT 334.150 1595.720 336.530 1596.370 ;
        RECT 337.370 1595.720 339.750 1596.370 ;
        RECT 340.590 1595.720 343.430 1596.370 ;
        RECT 344.270 1595.720 346.650 1596.370 ;
        RECT 347.490 1595.720 349.870 1596.370 ;
        RECT 350.710 1595.720 353.550 1596.370 ;
        RECT 354.390 1595.720 356.770 1596.370 ;
        RECT 357.610 1595.720 360.450 1596.370 ;
        RECT 361.290 1595.720 363.670 1596.370 ;
        RECT 364.510 1595.720 366.890 1596.370 ;
        RECT 367.730 1595.720 370.570 1596.370 ;
        RECT 371.410 1595.720 373.790 1596.370 ;
        RECT 374.630 1595.720 377.010 1596.370 ;
        RECT 377.850 1595.720 380.690 1596.370 ;
        RECT 381.530 1595.720 383.910 1596.370 ;
        RECT 384.750 1595.720 387.590 1596.370 ;
        RECT 388.430 1595.720 390.810 1596.370 ;
        RECT 391.650 1595.720 394.030 1596.370 ;
        RECT 394.870 1595.720 397.710 1596.370 ;
        RECT 398.550 1595.720 400.930 1596.370 ;
        RECT 401.770 1595.720 404.150 1596.370 ;
        RECT 404.990 1595.720 407.830 1596.370 ;
        RECT 408.670 1595.720 411.050 1596.370 ;
        RECT 411.890 1595.720 414.270 1596.370 ;
        RECT 415.110 1595.720 417.950 1596.370 ;
        RECT 418.790 1595.720 421.170 1596.370 ;
        RECT 422.010 1595.720 424.850 1596.370 ;
        RECT 425.690 1595.720 428.070 1596.370 ;
        RECT 428.910 1595.720 431.290 1596.370 ;
        RECT 432.130 1595.720 434.970 1596.370 ;
        RECT 435.810 1595.720 438.190 1596.370 ;
        RECT 439.030 1595.720 441.410 1596.370 ;
        RECT 442.250 1595.720 445.090 1596.370 ;
        RECT 445.930 1595.720 448.310 1596.370 ;
        RECT 449.150 1595.720 451.990 1596.370 ;
        RECT 452.830 1595.720 455.210 1596.370 ;
        RECT 456.050 1595.720 458.430 1596.370 ;
        RECT 459.270 1595.720 462.110 1596.370 ;
        RECT 462.950 1595.720 465.330 1596.370 ;
        RECT 466.170 1595.720 468.550 1596.370 ;
        RECT 469.390 1595.720 472.230 1596.370 ;
        RECT 473.070 1595.720 475.450 1596.370 ;
        RECT 476.290 1595.720 478.670 1596.370 ;
        RECT 479.510 1595.720 482.350 1596.370 ;
        RECT 483.190 1595.720 485.570 1596.370 ;
        RECT 486.410 1595.720 489.250 1596.370 ;
        RECT 490.090 1595.720 492.470 1596.370 ;
        RECT 493.310 1595.720 495.690 1596.370 ;
        RECT 496.530 1595.720 499.370 1596.370 ;
        RECT 500.210 1595.720 502.590 1596.370 ;
        RECT 503.430 1595.720 505.810 1596.370 ;
        RECT 506.650 1595.720 509.490 1596.370 ;
        RECT 510.330 1595.720 512.710 1596.370 ;
        RECT 513.550 1595.720 516.390 1596.370 ;
        RECT 517.230 1595.720 519.610 1596.370 ;
        RECT 520.450 1595.720 522.830 1596.370 ;
        RECT 523.670 1595.720 526.510 1596.370 ;
        RECT 527.350 1595.720 529.730 1596.370 ;
        RECT 530.570 1595.720 532.950 1596.370 ;
        RECT 533.790 1595.720 536.630 1596.370 ;
        RECT 537.470 1595.720 539.850 1596.370 ;
        RECT 540.690 1595.720 543.070 1596.370 ;
        RECT 543.910 1595.720 546.750 1596.370 ;
        RECT 547.590 1595.720 549.970 1596.370 ;
        RECT 550.810 1595.720 553.650 1596.370 ;
        RECT 554.490 1595.720 556.870 1596.370 ;
        RECT 557.710 1595.720 560.090 1596.370 ;
        RECT 560.930 1595.720 563.770 1596.370 ;
        RECT 564.610 1595.720 566.990 1596.370 ;
        RECT 567.830 1595.720 570.210 1596.370 ;
        RECT 571.050 1595.720 573.890 1596.370 ;
        RECT 574.730 1595.720 577.110 1596.370 ;
        RECT 577.950 1595.720 580.790 1596.370 ;
        RECT 581.630 1595.720 584.010 1596.370 ;
        RECT 584.850 1595.720 587.230 1596.370 ;
        RECT 588.070 1595.720 590.910 1596.370 ;
        RECT 591.750 1595.720 594.130 1596.370 ;
        RECT 594.970 1595.720 597.350 1596.370 ;
        RECT 598.190 1595.720 601.030 1596.370 ;
        RECT 601.870 1595.720 604.250 1596.370 ;
        RECT 605.090 1595.720 607.470 1596.370 ;
        RECT 608.310 1595.720 611.150 1596.370 ;
        RECT 611.990 1595.720 614.370 1596.370 ;
        RECT 615.210 1595.720 618.050 1596.370 ;
        RECT 618.890 1595.720 621.270 1596.370 ;
        RECT 622.110 1595.720 624.490 1596.370 ;
        RECT 625.330 1595.720 628.170 1596.370 ;
        RECT 629.010 1595.720 631.390 1596.370 ;
        RECT 632.230 1595.720 634.610 1596.370 ;
        RECT 635.450 1595.720 638.290 1596.370 ;
        RECT 639.130 1595.720 641.510 1596.370 ;
        RECT 642.350 1595.720 645.190 1596.370 ;
        RECT 646.030 1595.720 648.410 1596.370 ;
        RECT 649.250 1595.720 651.630 1596.370 ;
        RECT 652.470 1595.720 655.310 1596.370 ;
        RECT 656.150 1595.720 658.530 1596.370 ;
        RECT 659.370 1595.720 661.750 1596.370 ;
        RECT 662.590 1595.720 665.430 1596.370 ;
        RECT 666.270 1595.720 668.650 1596.370 ;
        RECT 669.490 1595.720 671.870 1596.370 ;
        RECT 672.710 1595.720 675.550 1596.370 ;
        RECT 676.390 1595.720 678.770 1596.370 ;
        RECT 679.610 1595.720 682.450 1596.370 ;
        RECT 683.290 1595.720 685.670 1596.370 ;
        RECT 686.510 1595.720 688.890 1596.370 ;
        RECT 689.730 1595.720 692.570 1596.370 ;
        RECT 693.410 1595.720 695.790 1596.370 ;
        RECT 696.630 1595.720 699.010 1596.370 ;
        RECT 699.850 1595.720 702.690 1596.370 ;
        RECT 703.530 1595.720 705.910 1596.370 ;
        RECT 706.750 1595.720 709.590 1596.370 ;
        RECT 710.430 1595.720 712.810 1596.370 ;
        RECT 713.650 1595.720 716.030 1596.370 ;
        RECT 716.870 1595.720 719.710 1596.370 ;
        RECT 720.550 1595.720 722.930 1596.370 ;
        RECT 723.770 1595.720 726.150 1596.370 ;
        RECT 726.990 1595.720 729.830 1596.370 ;
        RECT 730.670 1595.720 733.050 1596.370 ;
        RECT 733.890 1595.720 736.270 1596.370 ;
        RECT 737.110 1595.720 739.950 1596.370 ;
        RECT 740.790 1595.720 743.170 1596.370 ;
        RECT 744.010 1595.720 746.850 1596.370 ;
        RECT 747.690 1595.720 750.070 1596.370 ;
        RECT 750.910 1595.720 753.290 1596.370 ;
        RECT 754.130 1595.720 756.970 1596.370 ;
        RECT 757.810 1595.720 760.190 1596.370 ;
        RECT 761.030 1595.720 763.410 1596.370 ;
        RECT 764.250 1595.720 767.090 1596.370 ;
        RECT 767.930 1595.720 770.310 1596.370 ;
        RECT 771.150 1595.720 773.990 1596.370 ;
        RECT 774.830 1595.720 777.210 1596.370 ;
        RECT 778.050 1595.720 780.430 1596.370 ;
        RECT 781.270 1595.720 784.110 1596.370 ;
        RECT 784.950 1595.720 787.330 1596.370 ;
        RECT 788.170 1595.720 790.550 1596.370 ;
        RECT 791.390 1595.720 794.230 1596.370 ;
        RECT 0.100 4.280 794.780 1595.720 ;
        RECT 0.100 3.670 1.190 4.280 ;
        RECT 2.030 3.670 4.410 4.280 ;
        RECT 5.250 3.670 7.630 4.280 ;
        RECT 8.470 3.670 10.850 4.280 ;
        RECT 11.690 3.670 14.530 4.280 ;
        RECT 15.370 3.670 17.750 4.280 ;
        RECT 18.590 3.670 20.970 4.280 ;
        RECT 21.810 3.670 24.650 4.280 ;
        RECT 25.490 3.670 27.870 4.280 ;
        RECT 28.710 3.670 31.090 4.280 ;
        RECT 31.930 3.670 34.770 4.280 ;
        RECT 35.610 3.670 37.990 4.280 ;
        RECT 38.830 3.670 41.210 4.280 ;
        RECT 42.050 3.670 44.430 4.280 ;
        RECT 45.270 3.670 48.110 4.280 ;
        RECT 48.950 3.670 51.330 4.280 ;
        RECT 52.170 3.670 54.550 4.280 ;
        RECT 55.390 3.670 58.230 4.280 ;
        RECT 59.070 3.670 61.450 4.280 ;
        RECT 62.290 3.670 64.670 4.280 ;
        RECT 65.510 3.670 68.350 4.280 ;
        RECT 69.190 3.670 71.570 4.280 ;
        RECT 72.410 3.670 74.790 4.280 ;
        RECT 75.630 3.670 78.470 4.280 ;
        RECT 79.310 3.670 81.690 4.280 ;
        RECT 82.530 3.670 84.910 4.280 ;
        RECT 85.750 3.670 88.130 4.280 ;
        RECT 88.970 3.670 91.810 4.280 ;
        RECT 92.650 3.670 95.030 4.280 ;
        RECT 95.870 3.670 98.250 4.280 ;
        RECT 99.090 3.670 101.930 4.280 ;
        RECT 102.770 3.670 105.150 4.280 ;
        RECT 105.990 3.670 108.370 4.280 ;
        RECT 109.210 3.670 112.050 4.280 ;
        RECT 112.890 3.670 115.270 4.280 ;
        RECT 116.110 3.670 118.490 4.280 ;
        RECT 119.330 3.670 122.170 4.280 ;
        RECT 123.010 3.670 125.390 4.280 ;
        RECT 126.230 3.670 128.610 4.280 ;
        RECT 129.450 3.670 131.830 4.280 ;
        RECT 132.670 3.670 135.510 4.280 ;
        RECT 136.350 3.670 138.730 4.280 ;
        RECT 139.570 3.670 141.950 4.280 ;
        RECT 142.790 3.670 145.630 4.280 ;
        RECT 146.470 3.670 148.850 4.280 ;
        RECT 149.690 3.670 152.070 4.280 ;
        RECT 152.910 3.670 155.750 4.280 ;
        RECT 156.590 3.670 158.970 4.280 ;
        RECT 159.810 3.670 162.190 4.280 ;
        RECT 163.030 3.670 165.870 4.280 ;
        RECT 166.710 3.670 169.090 4.280 ;
        RECT 169.930 3.670 172.310 4.280 ;
        RECT 173.150 3.670 175.530 4.280 ;
        RECT 176.370 3.670 179.210 4.280 ;
        RECT 180.050 3.670 182.430 4.280 ;
        RECT 183.270 3.670 185.650 4.280 ;
        RECT 186.490 3.670 189.330 4.280 ;
        RECT 190.170 3.670 192.550 4.280 ;
        RECT 193.390 3.670 195.770 4.280 ;
        RECT 196.610 3.670 199.450 4.280 ;
        RECT 200.290 3.670 202.670 4.280 ;
        RECT 203.510 3.670 205.890 4.280 ;
        RECT 206.730 3.670 209.570 4.280 ;
        RECT 210.410 3.670 212.790 4.280 ;
        RECT 213.630 3.670 216.010 4.280 ;
        RECT 216.850 3.670 219.230 4.280 ;
        RECT 220.070 3.670 222.910 4.280 ;
        RECT 223.750 3.670 226.130 4.280 ;
        RECT 226.970 3.670 229.350 4.280 ;
        RECT 230.190 3.670 233.030 4.280 ;
        RECT 233.870 3.670 236.250 4.280 ;
        RECT 237.090 3.670 239.470 4.280 ;
        RECT 240.310 3.670 243.150 4.280 ;
        RECT 243.990 3.670 246.370 4.280 ;
        RECT 247.210 3.670 249.590 4.280 ;
        RECT 250.430 3.670 253.270 4.280 ;
        RECT 254.110 3.670 256.490 4.280 ;
        RECT 257.330 3.670 259.710 4.280 ;
        RECT 260.550 3.670 262.930 4.280 ;
        RECT 263.770 3.670 266.610 4.280 ;
        RECT 267.450 3.670 269.830 4.280 ;
        RECT 270.670 3.670 273.050 4.280 ;
        RECT 273.890 3.670 276.730 4.280 ;
        RECT 277.570 3.670 279.950 4.280 ;
        RECT 280.790 3.670 283.170 4.280 ;
        RECT 284.010 3.670 286.850 4.280 ;
        RECT 287.690 3.670 290.070 4.280 ;
        RECT 290.910 3.670 293.290 4.280 ;
        RECT 294.130 3.670 296.510 4.280 ;
        RECT 297.350 3.670 300.190 4.280 ;
        RECT 301.030 3.670 303.410 4.280 ;
        RECT 304.250 3.670 306.630 4.280 ;
        RECT 307.470 3.670 310.310 4.280 ;
        RECT 311.150 3.670 313.530 4.280 ;
        RECT 314.370 3.670 316.750 4.280 ;
        RECT 317.590 3.670 320.430 4.280 ;
        RECT 321.270 3.670 323.650 4.280 ;
        RECT 324.490 3.670 326.870 4.280 ;
        RECT 327.710 3.670 330.550 4.280 ;
        RECT 331.390 3.670 333.770 4.280 ;
        RECT 334.610 3.670 336.990 4.280 ;
        RECT 337.830 3.670 340.210 4.280 ;
        RECT 341.050 3.670 343.890 4.280 ;
        RECT 344.730 3.670 347.110 4.280 ;
        RECT 347.950 3.670 350.330 4.280 ;
        RECT 351.170 3.670 354.010 4.280 ;
        RECT 354.850 3.670 357.230 4.280 ;
        RECT 358.070 3.670 360.450 4.280 ;
        RECT 361.290 3.670 364.130 4.280 ;
        RECT 364.970 3.670 367.350 4.280 ;
        RECT 368.190 3.670 370.570 4.280 ;
        RECT 371.410 3.670 374.250 4.280 ;
        RECT 375.090 3.670 377.470 4.280 ;
        RECT 378.310 3.670 380.690 4.280 ;
        RECT 381.530 3.670 383.910 4.280 ;
        RECT 384.750 3.670 387.590 4.280 ;
        RECT 388.430 3.670 390.810 4.280 ;
        RECT 391.650 3.670 394.030 4.280 ;
        RECT 394.870 3.670 397.710 4.280 ;
        RECT 398.550 3.670 400.930 4.280 ;
        RECT 401.770 3.670 404.150 4.280 ;
        RECT 404.990 3.670 407.830 4.280 ;
        RECT 408.670 3.670 411.050 4.280 ;
        RECT 411.890 3.670 414.270 4.280 ;
        RECT 415.110 3.670 417.950 4.280 ;
        RECT 418.790 3.670 421.170 4.280 ;
        RECT 422.010 3.670 424.390 4.280 ;
        RECT 425.230 3.670 427.610 4.280 ;
        RECT 428.450 3.670 431.290 4.280 ;
        RECT 432.130 3.670 434.510 4.280 ;
        RECT 435.350 3.670 437.730 4.280 ;
        RECT 438.570 3.670 441.410 4.280 ;
        RECT 442.250 3.670 444.630 4.280 ;
        RECT 445.470 3.670 447.850 4.280 ;
        RECT 448.690 3.670 451.530 4.280 ;
        RECT 452.370 3.670 454.750 4.280 ;
        RECT 455.590 3.670 457.970 4.280 ;
        RECT 458.810 3.670 461.650 4.280 ;
        RECT 462.490 3.670 464.870 4.280 ;
        RECT 465.710 3.670 468.090 4.280 ;
        RECT 468.930 3.670 471.310 4.280 ;
        RECT 472.150 3.670 474.990 4.280 ;
        RECT 475.830 3.670 478.210 4.280 ;
        RECT 479.050 3.670 481.430 4.280 ;
        RECT 482.270 3.670 485.110 4.280 ;
        RECT 485.950 3.670 488.330 4.280 ;
        RECT 489.170 3.670 491.550 4.280 ;
        RECT 492.390 3.670 495.230 4.280 ;
        RECT 496.070 3.670 498.450 4.280 ;
        RECT 499.290 3.670 501.670 4.280 ;
        RECT 502.510 3.670 505.350 4.280 ;
        RECT 506.190 3.670 508.570 4.280 ;
        RECT 509.410 3.670 511.790 4.280 ;
        RECT 512.630 3.670 515.010 4.280 ;
        RECT 515.850 3.670 518.690 4.280 ;
        RECT 519.530 3.670 521.910 4.280 ;
        RECT 522.750 3.670 525.130 4.280 ;
        RECT 525.970 3.670 528.810 4.280 ;
        RECT 529.650 3.670 532.030 4.280 ;
        RECT 532.870 3.670 535.250 4.280 ;
        RECT 536.090 3.670 538.930 4.280 ;
        RECT 539.770 3.670 542.150 4.280 ;
        RECT 542.990 3.670 545.370 4.280 ;
        RECT 546.210 3.670 548.590 4.280 ;
        RECT 549.430 3.670 552.270 4.280 ;
        RECT 553.110 3.670 555.490 4.280 ;
        RECT 556.330 3.670 558.710 4.280 ;
        RECT 559.550 3.670 562.390 4.280 ;
        RECT 563.230 3.670 565.610 4.280 ;
        RECT 566.450 3.670 568.830 4.280 ;
        RECT 569.670 3.670 572.510 4.280 ;
        RECT 573.350 3.670 575.730 4.280 ;
        RECT 576.570 3.670 578.950 4.280 ;
        RECT 579.790 3.670 582.630 4.280 ;
        RECT 583.470 3.670 585.850 4.280 ;
        RECT 586.690 3.670 589.070 4.280 ;
        RECT 589.910 3.670 592.290 4.280 ;
        RECT 593.130 3.670 595.970 4.280 ;
        RECT 596.810 3.670 599.190 4.280 ;
        RECT 600.030 3.670 602.410 4.280 ;
        RECT 603.250 3.670 606.090 4.280 ;
        RECT 606.930 3.670 609.310 4.280 ;
        RECT 610.150 3.670 612.530 4.280 ;
        RECT 613.370 3.670 616.210 4.280 ;
        RECT 617.050 3.670 619.430 4.280 ;
        RECT 620.270 3.670 622.650 4.280 ;
        RECT 623.490 3.670 626.330 4.280 ;
        RECT 627.170 3.670 629.550 4.280 ;
        RECT 630.390 3.670 632.770 4.280 ;
        RECT 633.610 3.670 635.990 4.280 ;
        RECT 636.830 3.670 639.670 4.280 ;
        RECT 640.510 3.670 642.890 4.280 ;
        RECT 643.730 3.670 646.110 4.280 ;
        RECT 646.950 3.670 649.790 4.280 ;
        RECT 650.630 3.670 653.010 4.280 ;
        RECT 653.850 3.670 656.230 4.280 ;
        RECT 657.070 3.670 659.910 4.280 ;
        RECT 660.750 3.670 663.130 4.280 ;
        RECT 663.970 3.670 666.350 4.280 ;
        RECT 667.190 3.670 670.030 4.280 ;
        RECT 670.870 3.670 673.250 4.280 ;
        RECT 674.090 3.670 676.470 4.280 ;
        RECT 677.310 3.670 679.690 4.280 ;
        RECT 680.530 3.670 683.370 4.280 ;
        RECT 684.210 3.670 686.590 4.280 ;
        RECT 687.430 3.670 689.810 4.280 ;
        RECT 690.650 3.670 693.490 4.280 ;
        RECT 694.330 3.670 696.710 4.280 ;
        RECT 697.550 3.670 699.930 4.280 ;
        RECT 700.770 3.670 703.610 4.280 ;
        RECT 704.450 3.670 706.830 4.280 ;
        RECT 707.670 3.670 710.050 4.280 ;
        RECT 710.890 3.670 713.730 4.280 ;
        RECT 714.570 3.670 716.950 4.280 ;
        RECT 717.790 3.670 720.170 4.280 ;
        RECT 721.010 3.670 723.390 4.280 ;
        RECT 724.230 3.670 727.070 4.280 ;
        RECT 727.910 3.670 730.290 4.280 ;
        RECT 731.130 3.670 733.510 4.280 ;
        RECT 734.350 3.670 737.190 4.280 ;
        RECT 738.030 3.670 740.410 4.280 ;
        RECT 741.250 3.670 743.630 4.280 ;
        RECT 744.470 3.670 747.310 4.280 ;
        RECT 748.150 3.670 750.530 4.280 ;
        RECT 751.370 3.670 753.750 4.280 ;
        RECT 754.590 3.670 757.430 4.280 ;
        RECT 758.270 3.670 760.650 4.280 ;
        RECT 761.490 3.670 763.870 4.280 ;
        RECT 764.710 3.670 767.090 4.280 ;
        RECT 767.930 3.670 770.770 4.280 ;
        RECT 771.610 3.670 773.990 4.280 ;
        RECT 774.830 3.670 777.210 4.280 ;
        RECT 778.050 3.670 780.890 4.280 ;
        RECT 781.730 3.670 784.110 4.280 ;
        RECT 784.950 3.670 787.330 4.280 ;
        RECT 788.170 3.670 791.010 4.280 ;
        RECT 791.850 3.670 794.230 4.280 ;
      LAYER met3 ;
        RECT 4.000 1580.000 796.000 1588.645 ;
        RECT 4.400 1578.600 796.000 1580.000 ;
        RECT 4.000 1577.960 796.000 1578.600 ;
        RECT 4.000 1576.560 795.600 1577.960 ;
        RECT 4.000 1565.720 796.000 1576.560 ;
        RECT 4.400 1564.320 796.000 1565.720 ;
        RECT 4.000 1563.000 796.000 1564.320 ;
        RECT 4.000 1561.600 795.600 1563.000 ;
        RECT 4.000 1552.120 796.000 1561.600 ;
        RECT 4.400 1550.720 796.000 1552.120 ;
        RECT 4.000 1548.040 796.000 1550.720 ;
        RECT 4.000 1546.640 795.600 1548.040 ;
        RECT 4.000 1537.840 796.000 1546.640 ;
        RECT 4.400 1536.440 796.000 1537.840 ;
        RECT 4.000 1533.080 796.000 1536.440 ;
        RECT 4.000 1531.680 795.600 1533.080 ;
        RECT 4.000 1524.240 796.000 1531.680 ;
        RECT 4.400 1522.840 796.000 1524.240 ;
        RECT 4.000 1518.120 796.000 1522.840 ;
        RECT 4.000 1516.720 795.600 1518.120 ;
        RECT 4.000 1509.960 796.000 1516.720 ;
        RECT 4.400 1508.560 796.000 1509.960 ;
        RECT 4.000 1503.160 796.000 1508.560 ;
        RECT 4.000 1501.760 795.600 1503.160 ;
        RECT 4.000 1496.360 796.000 1501.760 ;
        RECT 4.400 1494.960 796.000 1496.360 ;
        RECT 4.000 1488.200 796.000 1494.960 ;
        RECT 4.000 1486.800 795.600 1488.200 ;
        RECT 4.000 1482.080 796.000 1486.800 ;
        RECT 4.400 1480.680 796.000 1482.080 ;
        RECT 4.000 1473.240 796.000 1480.680 ;
        RECT 4.000 1471.840 795.600 1473.240 ;
        RECT 4.000 1468.480 796.000 1471.840 ;
        RECT 4.400 1467.080 796.000 1468.480 ;
        RECT 4.000 1458.280 796.000 1467.080 ;
        RECT 4.000 1456.880 795.600 1458.280 ;
        RECT 4.000 1454.200 796.000 1456.880 ;
        RECT 4.400 1452.800 796.000 1454.200 ;
        RECT 4.000 1443.320 796.000 1452.800 ;
        RECT 4.000 1441.920 795.600 1443.320 ;
        RECT 4.000 1440.600 796.000 1441.920 ;
        RECT 4.400 1439.200 796.000 1440.600 ;
        RECT 4.000 1428.360 796.000 1439.200 ;
        RECT 4.000 1427.000 795.600 1428.360 ;
        RECT 4.400 1426.960 795.600 1427.000 ;
        RECT 4.400 1425.600 796.000 1426.960 ;
        RECT 4.000 1413.400 796.000 1425.600 ;
        RECT 4.000 1412.720 795.600 1413.400 ;
        RECT 4.400 1412.000 795.600 1412.720 ;
        RECT 4.400 1411.320 796.000 1412.000 ;
        RECT 4.000 1399.120 796.000 1411.320 ;
        RECT 4.400 1398.440 796.000 1399.120 ;
        RECT 4.400 1397.720 795.600 1398.440 ;
        RECT 4.000 1397.040 795.600 1397.720 ;
        RECT 4.000 1384.840 796.000 1397.040 ;
        RECT 4.400 1383.480 796.000 1384.840 ;
        RECT 4.400 1383.440 795.600 1383.480 ;
        RECT 4.000 1382.080 795.600 1383.440 ;
        RECT 4.000 1371.240 796.000 1382.080 ;
        RECT 4.400 1369.840 796.000 1371.240 ;
        RECT 4.000 1368.520 796.000 1369.840 ;
        RECT 4.000 1367.120 795.600 1368.520 ;
        RECT 4.000 1356.960 796.000 1367.120 ;
        RECT 4.400 1355.560 796.000 1356.960 ;
        RECT 4.000 1353.560 796.000 1355.560 ;
        RECT 4.000 1352.160 795.600 1353.560 ;
        RECT 4.000 1343.360 796.000 1352.160 ;
        RECT 4.400 1341.960 796.000 1343.360 ;
        RECT 4.000 1338.600 796.000 1341.960 ;
        RECT 4.000 1337.200 795.600 1338.600 ;
        RECT 4.000 1329.080 796.000 1337.200 ;
        RECT 4.400 1327.680 796.000 1329.080 ;
        RECT 4.000 1323.640 796.000 1327.680 ;
        RECT 4.000 1322.240 795.600 1323.640 ;
        RECT 4.000 1315.480 796.000 1322.240 ;
        RECT 4.400 1314.080 796.000 1315.480 ;
        RECT 4.000 1308.680 796.000 1314.080 ;
        RECT 4.000 1307.280 795.600 1308.680 ;
        RECT 4.000 1301.200 796.000 1307.280 ;
        RECT 4.400 1299.800 796.000 1301.200 ;
        RECT 4.000 1293.720 796.000 1299.800 ;
        RECT 4.000 1292.320 795.600 1293.720 ;
        RECT 4.000 1287.600 796.000 1292.320 ;
        RECT 4.400 1286.200 796.000 1287.600 ;
        RECT 4.000 1278.760 796.000 1286.200 ;
        RECT 4.000 1277.360 795.600 1278.760 ;
        RECT 4.000 1273.320 796.000 1277.360 ;
        RECT 4.400 1271.920 796.000 1273.320 ;
        RECT 4.000 1263.800 796.000 1271.920 ;
        RECT 4.000 1262.400 795.600 1263.800 ;
        RECT 4.000 1259.720 796.000 1262.400 ;
        RECT 4.400 1258.320 796.000 1259.720 ;
        RECT 4.000 1248.840 796.000 1258.320 ;
        RECT 4.000 1247.440 795.600 1248.840 ;
        RECT 4.000 1246.120 796.000 1247.440 ;
        RECT 4.400 1244.720 796.000 1246.120 ;
        RECT 4.000 1233.880 796.000 1244.720 ;
        RECT 4.000 1232.480 795.600 1233.880 ;
        RECT 4.000 1231.840 796.000 1232.480 ;
        RECT 4.400 1230.440 796.000 1231.840 ;
        RECT 4.000 1218.920 796.000 1230.440 ;
        RECT 4.000 1218.240 795.600 1218.920 ;
        RECT 4.400 1217.520 795.600 1218.240 ;
        RECT 4.400 1216.840 796.000 1217.520 ;
        RECT 4.000 1203.960 796.000 1216.840 ;
        RECT 4.400 1202.560 795.600 1203.960 ;
        RECT 4.000 1190.360 796.000 1202.560 ;
        RECT 4.400 1189.000 796.000 1190.360 ;
        RECT 4.400 1188.960 795.600 1189.000 ;
        RECT 4.000 1187.600 795.600 1188.960 ;
        RECT 4.000 1176.080 796.000 1187.600 ;
        RECT 4.400 1174.680 796.000 1176.080 ;
        RECT 4.000 1174.040 796.000 1174.680 ;
        RECT 4.000 1172.640 795.600 1174.040 ;
        RECT 4.000 1162.480 796.000 1172.640 ;
        RECT 4.400 1161.080 796.000 1162.480 ;
        RECT 4.000 1159.080 796.000 1161.080 ;
        RECT 4.000 1157.680 795.600 1159.080 ;
        RECT 4.000 1148.200 796.000 1157.680 ;
        RECT 4.400 1146.800 796.000 1148.200 ;
        RECT 4.000 1144.120 796.000 1146.800 ;
        RECT 4.000 1142.720 795.600 1144.120 ;
        RECT 4.000 1134.600 796.000 1142.720 ;
        RECT 4.400 1133.200 796.000 1134.600 ;
        RECT 4.000 1129.160 796.000 1133.200 ;
        RECT 4.000 1127.760 795.600 1129.160 ;
        RECT 4.000 1120.320 796.000 1127.760 ;
        RECT 4.400 1118.920 796.000 1120.320 ;
        RECT 4.000 1114.200 796.000 1118.920 ;
        RECT 4.000 1112.800 795.600 1114.200 ;
        RECT 4.000 1106.720 796.000 1112.800 ;
        RECT 4.400 1105.320 796.000 1106.720 ;
        RECT 4.000 1099.240 796.000 1105.320 ;
        RECT 4.000 1097.840 795.600 1099.240 ;
        RECT 4.000 1092.440 796.000 1097.840 ;
        RECT 4.400 1091.040 796.000 1092.440 ;
        RECT 4.000 1084.280 796.000 1091.040 ;
        RECT 4.000 1082.880 795.600 1084.280 ;
        RECT 4.000 1078.840 796.000 1082.880 ;
        RECT 4.400 1077.440 796.000 1078.840 ;
        RECT 4.000 1069.320 796.000 1077.440 ;
        RECT 4.000 1067.920 795.600 1069.320 ;
        RECT 4.000 1065.240 796.000 1067.920 ;
        RECT 4.400 1063.840 796.000 1065.240 ;
        RECT 4.000 1054.360 796.000 1063.840 ;
        RECT 4.000 1052.960 795.600 1054.360 ;
        RECT 4.000 1050.960 796.000 1052.960 ;
        RECT 4.400 1049.560 796.000 1050.960 ;
        RECT 4.000 1039.400 796.000 1049.560 ;
        RECT 4.000 1038.000 795.600 1039.400 ;
        RECT 4.000 1037.360 796.000 1038.000 ;
        RECT 4.400 1035.960 796.000 1037.360 ;
        RECT 4.000 1024.440 796.000 1035.960 ;
        RECT 4.000 1023.080 795.600 1024.440 ;
        RECT 4.400 1023.040 795.600 1023.080 ;
        RECT 4.400 1021.680 796.000 1023.040 ;
        RECT 4.000 1009.480 796.000 1021.680 ;
        RECT 4.400 1008.080 795.600 1009.480 ;
        RECT 4.000 995.200 796.000 1008.080 ;
        RECT 4.400 994.520 796.000 995.200 ;
        RECT 4.400 993.800 795.600 994.520 ;
        RECT 4.000 993.120 795.600 993.800 ;
        RECT 4.000 981.600 796.000 993.120 ;
        RECT 4.400 980.200 796.000 981.600 ;
        RECT 4.000 979.560 796.000 980.200 ;
        RECT 4.000 978.160 795.600 979.560 ;
        RECT 4.000 967.320 796.000 978.160 ;
        RECT 4.400 965.920 796.000 967.320 ;
        RECT 4.000 964.600 796.000 965.920 ;
        RECT 4.000 963.200 795.600 964.600 ;
        RECT 4.000 953.720 796.000 963.200 ;
        RECT 4.400 952.320 796.000 953.720 ;
        RECT 4.000 949.640 796.000 952.320 ;
        RECT 4.000 948.240 795.600 949.640 ;
        RECT 4.000 939.440 796.000 948.240 ;
        RECT 4.400 938.040 796.000 939.440 ;
        RECT 4.000 934.680 796.000 938.040 ;
        RECT 4.000 933.280 795.600 934.680 ;
        RECT 4.000 925.840 796.000 933.280 ;
        RECT 4.400 924.440 796.000 925.840 ;
        RECT 4.000 919.720 796.000 924.440 ;
        RECT 4.000 918.320 795.600 919.720 ;
        RECT 4.000 911.560 796.000 918.320 ;
        RECT 4.400 910.160 796.000 911.560 ;
        RECT 4.000 904.760 796.000 910.160 ;
        RECT 4.000 903.360 795.600 904.760 ;
        RECT 4.000 897.960 796.000 903.360 ;
        RECT 4.400 896.560 796.000 897.960 ;
        RECT 4.000 889.800 796.000 896.560 ;
        RECT 4.000 888.400 795.600 889.800 ;
        RECT 4.000 884.360 796.000 888.400 ;
        RECT 4.400 882.960 796.000 884.360 ;
        RECT 4.000 874.840 796.000 882.960 ;
        RECT 4.000 873.440 795.600 874.840 ;
        RECT 4.000 870.080 796.000 873.440 ;
        RECT 4.400 868.680 796.000 870.080 ;
        RECT 4.000 859.880 796.000 868.680 ;
        RECT 4.000 858.480 795.600 859.880 ;
        RECT 4.000 856.480 796.000 858.480 ;
        RECT 4.400 855.080 796.000 856.480 ;
        RECT 4.000 844.920 796.000 855.080 ;
        RECT 4.000 843.520 795.600 844.920 ;
        RECT 4.000 842.200 796.000 843.520 ;
        RECT 4.400 840.800 796.000 842.200 ;
        RECT 4.000 829.960 796.000 840.800 ;
        RECT 4.000 828.600 795.600 829.960 ;
        RECT 4.400 828.560 795.600 828.600 ;
        RECT 4.400 827.200 796.000 828.560 ;
        RECT 4.000 815.000 796.000 827.200 ;
        RECT 4.000 814.320 795.600 815.000 ;
        RECT 4.400 813.600 795.600 814.320 ;
        RECT 4.400 812.920 796.000 813.600 ;
        RECT 4.000 800.720 796.000 812.920 ;
        RECT 4.400 800.040 796.000 800.720 ;
        RECT 4.400 799.320 795.600 800.040 ;
        RECT 4.000 798.640 795.600 799.320 ;
        RECT 4.000 786.440 796.000 798.640 ;
        RECT 4.400 785.080 796.000 786.440 ;
        RECT 4.400 785.040 795.600 785.080 ;
        RECT 4.000 783.680 795.600 785.040 ;
        RECT 4.000 772.840 796.000 783.680 ;
        RECT 4.400 771.440 796.000 772.840 ;
        RECT 4.000 770.120 796.000 771.440 ;
        RECT 4.000 768.720 795.600 770.120 ;
        RECT 4.000 758.560 796.000 768.720 ;
        RECT 4.400 757.160 796.000 758.560 ;
        RECT 4.000 755.160 796.000 757.160 ;
        RECT 4.000 753.760 795.600 755.160 ;
        RECT 4.000 744.960 796.000 753.760 ;
        RECT 4.400 743.560 796.000 744.960 ;
        RECT 4.000 740.200 796.000 743.560 ;
        RECT 4.000 738.800 795.600 740.200 ;
        RECT 4.000 730.680 796.000 738.800 ;
        RECT 4.400 729.280 796.000 730.680 ;
        RECT 4.000 725.240 796.000 729.280 ;
        RECT 4.000 723.840 795.600 725.240 ;
        RECT 4.000 717.080 796.000 723.840 ;
        RECT 4.400 715.680 796.000 717.080 ;
        RECT 4.000 710.280 796.000 715.680 ;
        RECT 4.000 708.880 795.600 710.280 ;
        RECT 4.000 703.480 796.000 708.880 ;
        RECT 4.400 702.080 796.000 703.480 ;
        RECT 4.000 695.320 796.000 702.080 ;
        RECT 4.000 693.920 795.600 695.320 ;
        RECT 4.000 689.200 796.000 693.920 ;
        RECT 4.400 687.800 796.000 689.200 ;
        RECT 4.000 680.360 796.000 687.800 ;
        RECT 4.000 678.960 795.600 680.360 ;
        RECT 4.000 675.600 796.000 678.960 ;
        RECT 4.400 674.200 796.000 675.600 ;
        RECT 4.000 665.400 796.000 674.200 ;
        RECT 4.000 664.000 795.600 665.400 ;
        RECT 4.000 661.320 796.000 664.000 ;
        RECT 4.400 659.920 796.000 661.320 ;
        RECT 4.000 650.440 796.000 659.920 ;
        RECT 4.000 649.040 795.600 650.440 ;
        RECT 4.000 647.720 796.000 649.040 ;
        RECT 4.400 646.320 796.000 647.720 ;
        RECT 4.000 635.480 796.000 646.320 ;
        RECT 4.000 634.080 795.600 635.480 ;
        RECT 4.000 633.440 796.000 634.080 ;
        RECT 4.400 632.040 796.000 633.440 ;
        RECT 4.000 620.520 796.000 632.040 ;
        RECT 4.000 619.840 795.600 620.520 ;
        RECT 4.400 619.120 795.600 619.840 ;
        RECT 4.400 618.440 796.000 619.120 ;
        RECT 4.000 605.560 796.000 618.440 ;
        RECT 4.400 604.160 795.600 605.560 ;
        RECT 4.000 591.960 796.000 604.160 ;
        RECT 4.400 590.600 796.000 591.960 ;
        RECT 4.400 590.560 795.600 590.600 ;
        RECT 4.000 589.200 795.600 590.560 ;
        RECT 4.000 577.680 796.000 589.200 ;
        RECT 4.400 576.280 796.000 577.680 ;
        RECT 4.000 575.640 796.000 576.280 ;
        RECT 4.000 574.240 795.600 575.640 ;
        RECT 4.000 564.080 796.000 574.240 ;
        RECT 4.400 562.680 796.000 564.080 ;
        RECT 4.000 560.680 796.000 562.680 ;
        RECT 4.000 559.280 795.600 560.680 ;
        RECT 4.000 549.800 796.000 559.280 ;
        RECT 4.400 548.400 796.000 549.800 ;
        RECT 4.000 545.720 796.000 548.400 ;
        RECT 4.000 544.320 795.600 545.720 ;
        RECT 4.000 536.200 796.000 544.320 ;
        RECT 4.400 534.800 796.000 536.200 ;
        RECT 4.000 530.760 796.000 534.800 ;
        RECT 4.000 529.360 795.600 530.760 ;
        RECT 4.000 522.600 796.000 529.360 ;
        RECT 4.400 521.200 796.000 522.600 ;
        RECT 4.000 515.800 796.000 521.200 ;
        RECT 4.000 514.400 795.600 515.800 ;
        RECT 4.000 508.320 796.000 514.400 ;
        RECT 4.400 506.920 796.000 508.320 ;
        RECT 4.000 500.840 796.000 506.920 ;
        RECT 4.000 499.440 795.600 500.840 ;
        RECT 4.000 494.720 796.000 499.440 ;
        RECT 4.400 493.320 796.000 494.720 ;
        RECT 4.000 485.880 796.000 493.320 ;
        RECT 4.000 484.480 795.600 485.880 ;
        RECT 4.000 480.440 796.000 484.480 ;
        RECT 4.400 479.040 796.000 480.440 ;
        RECT 4.000 470.920 796.000 479.040 ;
        RECT 4.000 469.520 795.600 470.920 ;
        RECT 4.000 466.840 796.000 469.520 ;
        RECT 4.400 465.440 796.000 466.840 ;
        RECT 4.000 455.960 796.000 465.440 ;
        RECT 4.000 454.560 795.600 455.960 ;
        RECT 4.000 452.560 796.000 454.560 ;
        RECT 4.400 451.160 796.000 452.560 ;
        RECT 4.000 441.000 796.000 451.160 ;
        RECT 4.000 439.600 795.600 441.000 ;
        RECT 4.000 438.960 796.000 439.600 ;
        RECT 4.400 437.560 796.000 438.960 ;
        RECT 4.000 426.040 796.000 437.560 ;
        RECT 4.000 424.680 795.600 426.040 ;
        RECT 4.400 424.640 795.600 424.680 ;
        RECT 4.400 423.280 796.000 424.640 ;
        RECT 4.000 411.080 796.000 423.280 ;
        RECT 4.400 409.680 795.600 411.080 ;
        RECT 4.000 396.800 796.000 409.680 ;
        RECT 4.400 396.120 796.000 396.800 ;
        RECT 4.400 395.400 795.600 396.120 ;
        RECT 4.000 394.720 795.600 395.400 ;
        RECT 4.000 383.200 796.000 394.720 ;
        RECT 4.400 381.800 796.000 383.200 ;
        RECT 4.000 381.160 796.000 381.800 ;
        RECT 4.000 379.760 795.600 381.160 ;
        RECT 4.000 368.920 796.000 379.760 ;
        RECT 4.400 367.520 796.000 368.920 ;
        RECT 4.000 366.200 796.000 367.520 ;
        RECT 4.000 364.800 795.600 366.200 ;
        RECT 4.000 355.320 796.000 364.800 ;
        RECT 4.400 353.920 796.000 355.320 ;
        RECT 4.000 351.240 796.000 353.920 ;
        RECT 4.000 349.840 795.600 351.240 ;
        RECT 4.000 341.720 796.000 349.840 ;
        RECT 4.400 340.320 796.000 341.720 ;
        RECT 4.000 336.280 796.000 340.320 ;
        RECT 4.000 334.880 795.600 336.280 ;
        RECT 4.000 327.440 796.000 334.880 ;
        RECT 4.400 326.040 796.000 327.440 ;
        RECT 4.000 321.320 796.000 326.040 ;
        RECT 4.000 319.920 795.600 321.320 ;
        RECT 4.000 313.840 796.000 319.920 ;
        RECT 4.400 312.440 796.000 313.840 ;
        RECT 4.000 306.360 796.000 312.440 ;
        RECT 4.000 304.960 795.600 306.360 ;
        RECT 4.000 299.560 796.000 304.960 ;
        RECT 4.400 298.160 796.000 299.560 ;
        RECT 4.000 291.400 796.000 298.160 ;
        RECT 4.000 290.000 795.600 291.400 ;
        RECT 4.000 285.960 796.000 290.000 ;
        RECT 4.400 284.560 796.000 285.960 ;
        RECT 4.000 276.440 796.000 284.560 ;
        RECT 4.000 275.040 795.600 276.440 ;
        RECT 4.000 271.680 796.000 275.040 ;
        RECT 4.400 270.280 796.000 271.680 ;
        RECT 4.000 261.480 796.000 270.280 ;
        RECT 4.000 260.080 795.600 261.480 ;
        RECT 4.000 258.080 796.000 260.080 ;
        RECT 4.400 256.680 796.000 258.080 ;
        RECT 4.000 246.520 796.000 256.680 ;
        RECT 4.000 245.120 795.600 246.520 ;
        RECT 4.000 243.800 796.000 245.120 ;
        RECT 4.400 242.400 796.000 243.800 ;
        RECT 4.000 231.560 796.000 242.400 ;
        RECT 4.000 230.200 795.600 231.560 ;
        RECT 4.400 230.160 795.600 230.200 ;
        RECT 4.400 228.800 796.000 230.160 ;
        RECT 4.000 216.600 796.000 228.800 ;
        RECT 4.000 215.920 795.600 216.600 ;
        RECT 4.400 215.200 795.600 215.920 ;
        RECT 4.400 214.520 796.000 215.200 ;
        RECT 4.000 202.320 796.000 214.520 ;
        RECT 4.400 201.640 796.000 202.320 ;
        RECT 4.400 200.920 795.600 201.640 ;
        RECT 4.000 200.240 795.600 200.920 ;
        RECT 4.000 188.040 796.000 200.240 ;
        RECT 4.400 186.680 796.000 188.040 ;
        RECT 4.400 186.640 795.600 186.680 ;
        RECT 4.000 185.280 795.600 186.640 ;
        RECT 4.000 174.440 796.000 185.280 ;
        RECT 4.400 173.040 796.000 174.440 ;
        RECT 4.000 171.720 796.000 173.040 ;
        RECT 4.000 170.320 795.600 171.720 ;
        RECT 4.000 160.840 796.000 170.320 ;
        RECT 4.400 159.440 796.000 160.840 ;
        RECT 4.000 156.760 796.000 159.440 ;
        RECT 4.000 155.360 795.600 156.760 ;
        RECT 4.000 146.560 796.000 155.360 ;
        RECT 4.400 145.160 796.000 146.560 ;
        RECT 4.000 141.800 796.000 145.160 ;
        RECT 4.000 140.400 795.600 141.800 ;
        RECT 4.000 132.960 796.000 140.400 ;
        RECT 4.400 131.560 796.000 132.960 ;
        RECT 4.000 126.840 796.000 131.560 ;
        RECT 4.000 125.440 795.600 126.840 ;
        RECT 4.000 118.680 796.000 125.440 ;
        RECT 4.400 117.280 796.000 118.680 ;
        RECT 4.000 111.880 796.000 117.280 ;
        RECT 4.000 110.480 795.600 111.880 ;
        RECT 4.000 105.080 796.000 110.480 ;
        RECT 4.400 103.680 796.000 105.080 ;
        RECT 4.000 96.920 796.000 103.680 ;
        RECT 4.000 95.520 795.600 96.920 ;
        RECT 4.000 90.800 796.000 95.520 ;
        RECT 4.400 89.400 796.000 90.800 ;
        RECT 4.000 81.960 796.000 89.400 ;
        RECT 4.000 80.560 795.600 81.960 ;
        RECT 4.000 77.200 796.000 80.560 ;
        RECT 4.400 75.800 796.000 77.200 ;
        RECT 4.000 67.000 796.000 75.800 ;
        RECT 4.000 65.600 795.600 67.000 ;
        RECT 4.000 62.920 796.000 65.600 ;
        RECT 4.400 61.520 796.000 62.920 ;
        RECT 4.000 52.040 796.000 61.520 ;
        RECT 4.000 50.640 795.600 52.040 ;
        RECT 4.000 49.320 796.000 50.640 ;
        RECT 4.400 47.920 796.000 49.320 ;
        RECT 4.000 37.080 796.000 47.920 ;
        RECT 4.000 35.680 795.600 37.080 ;
        RECT 4.000 35.040 796.000 35.680 ;
        RECT 4.400 33.640 796.000 35.040 ;
        RECT 4.000 22.120 796.000 33.640 ;
        RECT 4.000 21.440 795.600 22.120 ;
        RECT 4.400 20.720 795.600 21.440 ;
        RECT 4.400 20.040 796.000 20.720 ;
        RECT 4.000 7.840 796.000 20.040 ;
        RECT 4.400 6.975 795.600 7.840 ;
      LAYER met4 ;
        RECT 163.135 27.375 174.240 592.105 ;
        RECT 176.640 27.375 250.865 592.105 ;
  END
END user_proj_example
END LIBRARY

