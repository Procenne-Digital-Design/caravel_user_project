VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 1600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 836.440 800.000 837.040 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 635.840 800.000 636.440 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1596.000 193.570 1600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1596.000 251.530 1600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1596.000 309.490 1600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1020.040 800.000 1020.640 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 724.240 800.000 724.840 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 972.440 800.000 973.040 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 285.640 800.000 286.240 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 513.440 800.000 514.040 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 1596.000 731.310 1600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 425.040 800.000 425.640 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 95.240 800.000 95.840 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 1596.000 789.270 1600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 1596.000 71.210 1600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 299.240 800.000 299.840 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.040 4.000 1224.640 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 231.240 800.000 231.840 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 918.040 800.000 918.640 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 1596.000 96.970 1600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1530.040 4.000 1530.640 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1292.040 4.000 1292.640 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1596.000 39.010 1600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 1596.000 769.950 1600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 1596.000 660.470 1600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 1596.000 505.910 1600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1540.240 800.000 1540.840 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1370.240 800.000 1370.840 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1570.840 4.000 1571.440 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1424.640 800.000 1425.240 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1142.440 800.000 1143.040 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1591.240 4.000 1591.840 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1596.000 737.750 1600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 340.040 800.000 340.640 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1094.840 800.000 1095.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 1596.000 557.430 1600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.840 800.000 177.440 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 68.040 800.000 68.640 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 1596.000 493.030 1600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1451.840 800.000 1452.440 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 904.440 800.000 905.040 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.040 4.000 1496.640 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1567.440 800.000 1568.040 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 1596.000 277.290 1600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 758.240 800.000 758.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 102.040 800.000 102.640 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 744.640 800.000 745.240 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1553.840 800.000 1554.440 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1207.040 800.000 1207.640 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1574.240 800.000 1574.840 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1596.000 64.770 1600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 1596.000 245.090 1600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1081.240 800.000 1081.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1596.000 460.830 1600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 20.440 800.000 21.040 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 1596.000 795.710 1600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1458.640 800.000 1459.240 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 1596.000 270.850 1600.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 1596.000 563.870 1600.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 1596.000 264.410 1600.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 1596.000 206.450 1600.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1596.000 570.310 1600.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 88.440 800.000 89.040 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 1596.000 724.870 1600.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 843.240 800.000 843.840 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 622.240 800.000 622.840 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 486.240 800.000 486.840 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 608.640 800.000 609.240 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 1596.000 412.530 1600.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 1596.000 84.090 1600.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1596.000 167.810 1600.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1596.000 22.910 1600.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1054.040 800.000 1054.640 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 676.640 800.000 677.240 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 190.440 800.000 191.040 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 384.240 800.000 384.840 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 1596.000 348.130 1600.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 1596.000 750.630 1600.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 1596.000 187.130 1600.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1115.240 800.000 1115.840 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 999.640 800.000 1000.240 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1067.640 800.000 1068.240 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 649.440 800.000 650.040 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1200.240 800.000 1200.840 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1149.240 800.000 1149.840 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1596.000 480.150 1600.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1596.000 225.770 1600.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 1596.000 634.710 1600.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1213.840 800.000 1214.440 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 404.640 800.000 405.240 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 938.440 800.000 939.040 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 1596.000 576.750 1600.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 1596.000 290.170 1600.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 81.640 800.000 82.240 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1596.000 135.610 1600.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1499.440 800.000 1500.040 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 554.240 800.000 554.840 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1596.000 16.470 1600.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1596.000 531.670 1600.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1587.840 800.000 1588.440 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 1596.000 447.950 1600.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1596.000 174.250 1600.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 690.240 800.000 690.840 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 452.240 800.000 452.840 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1390.640 800.000 1391.240 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1241.040 800.000 1241.640 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1431.440 800.000 1432.040 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1596.000 161.370 1600.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1414.440 4.000 1415.040 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 506.640 800.000 507.240 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1278.440 4.000 1279.040 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 1596.000 406.090 1600.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1596.000 782.830 1600.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1596.000 386.770 1600.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 1596.000 393.210 1600.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1183.240 800.000 1183.840 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 360.440 800.000 361.040 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 1596.000 718.430 1600.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1336.240 800.000 1336.840 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 877.240 800.000 877.840 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 1596.000 699.110 1600.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1596.000 148.490 1600.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 809.240 800.000 809.840 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 778.640 800.000 779.240 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 663.040 800.000 663.640 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 897.640 800.000 898.240 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1596.000 467.270 1600.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1596.000 129.170 1600.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 1596.000 303.050 1600.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1596.000 154.930 1600.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1596.000 122.730 1600.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 353.640 800.000 354.240 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1383.840 800.000 1384.440 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 642.640 800.000 643.240 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1006.440 800.000 1007.040 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 1596.000 596.070 1600.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 1596.000 238.650 1600.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1596.000 673.350 1600.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 122.440 800.000 123.040 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1596.000 550.990 1600.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 1596.000 602.510 1600.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1596.000 776.390 1600.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 1596.000 435.070 1600.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 326.440 800.000 327.040 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 1596.000 679.790 1600.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 292.440 800.000 293.040 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 1596.000 711.990 1600.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 771.840 800.000 772.440 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1596.000 109.850 1600.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 952.040 800.000 952.640 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 945.240 800.000 945.840 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 244.840 800.000 245.440 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1445.040 800.000 1445.640 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1596.000 621.830 1600.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 1596.000 373.890 1600.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 108.840 800.000 109.440 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1596.000 45.450 1600.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 238.040 800.000 238.640 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1465.440 800.000 1466.040 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1533.440 800.000 1534.040 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 540.640 800.000 541.240 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 795.640 800.000 796.240 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1438.240 800.000 1438.840 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 418.240 800.000 418.840 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1596.000 200.010 1600.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 129.240 800.000 129.840 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 581.440 800.000 582.040 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1315.840 800.000 1316.440 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1169.640 800.000 1170.240 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 472.640 800.000 473.240 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 61.240 800.000 61.840 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1417.840 800.000 1418.440 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1322.640 800.000 1323.240 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1135.640 800.000 1136.240 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1411.040 800.000 1411.640 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 391.040 800.000 391.640 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 588.240 800.000 588.840 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.840 4.000 1469.440 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1190.040 800.000 1190.640 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1108.440 800.000 1109.040 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1596.000 544.550 1600.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 47.640 800.000 48.240 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1122.040 800.000 1122.640 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1060.840 800.000 1061.440 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1596.000 518.790 1600.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1047.240 800.000 1047.840 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 785.440 800.000 786.040 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1547.040 800.000 1547.640 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 601.840 800.000 602.440 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1176.440 800.000 1177.040 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1220.640 800.000 1221.240 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 438.640 800.000 439.240 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1596.000 692.670 1600.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1596.000 666.910 1600.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1584.440 4.000 1585.040 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 374.040 800.000 374.640 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1101.640 800.000 1102.240 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 731.040 800.000 731.640 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 1596.000 686.230 1600.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1404.240 800.000 1404.840 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 958.840 800.000 959.440 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.040 4.000 1598.640 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 816.040 800.000 816.640 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1485.840 800.000 1486.440 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 445.440 800.000 446.040 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.040 4.000 1207.640 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 1596.000 322.370 1600.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 788.840 800.000 789.440 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1596.000 315.930 1600.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 465.840 800.000 466.440 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 4.000 1251.840 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 911.240 800.000 911.840 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 697.040 800.000 697.640 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 986.040 800.000 986.640 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1596.000 26.130 1600.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1377.040 800.000 1377.640 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1281.840 800.000 1282.440 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 224.440 800.000 225.040 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 863.640 800.000 864.240 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 870.440 800.000 871.040 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 431.840 800.000 432.440 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 156.440 800.000 157.040 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1156.040 800.000 1156.640 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1186.640 4.000 1187.240 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1261.440 800.000 1262.040 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1026.840 800.000 1027.440 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 703.840 800.000 704.440 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 4.000 1245.040 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 411.440 800.000 412.040 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 533.840 800.000 534.440 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 656.240 800.000 656.840 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1088.040 800.000 1088.640 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1596.000 212.890 1600.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 346.840 800.000 347.440 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 615.440 800.000 616.040 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 1596.000 422.190 1600.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1237.640 4.000 1238.240 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1268.240 800.000 1268.840 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 629.040 800.000 629.640 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1596.000 77.650 1600.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1596.000 341.690 1600.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 377.440 800.000 378.040 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1288.640 800.000 1289.240 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 197.240 800.000 197.840 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1309.040 800.000 1309.640 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 459.040 800.000 459.640 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 765.040 800.000 765.640 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 115.640 800.000 116.240 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1596.000 525.230 1600.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 272.040 800.000 272.640 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 1596.000 647.590 1600.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 520.240 800.000 520.840 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 27.240 800.000 27.840 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1596.000 335.250 1600.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 183.640 800.000 184.240 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 312.840 800.000 313.440 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 1596.000 354.570 1600.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1596.000 615.390 1600.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 924.840 800.000 925.440 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 1596.000 328.810 1600.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1596.000 583.190 1600.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 669.840 800.000 670.440 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 1596.000 361.010 1600.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1275.040 800.000 1275.640 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 142.840 800.000 143.440 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END la_oenb[9]
  PIN sram_addr_a[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 1596.000 142.050 1600.000 ;
    END
  END sram_addr_a[0]
  PIN sram_addr_a[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END sram_addr_a[1]
  PIN sram_addr_a[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END sram_addr_a[2]
  PIN sram_addr_a[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1513.040 800.000 1513.640 ;
    END
  END sram_addr_a[3]
  PIN sram_addr_a[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 136.040 800.000 136.640 ;
    END
  END sram_addr_a[4]
  PIN sram_addr_a[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END sram_addr_a[5]
  PIN sram_addr_a[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END sram_addr_a[6]
  PIN sram_addr_a[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END sram_addr_a[7]
  PIN sram_addr_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END sram_addr_b[0]
  PIN sram_addr_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END sram_addr_b[1]
  PIN sram_addr_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1596.000 654.030 1600.000 ;
    END
  END sram_addr_b[2]
  PIN sram_addr_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1013.240 800.000 1013.840 ;
    END
  END sram_addr_b[3]
  PIN sram_addr_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 567.840 800.000 568.440 ;
    END
  END sram_addr_b[4]
  PIN sram_addr_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1247.840 800.000 1248.440 ;
    END
  END sram_addr_b[5]
  PIN sram_addr_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 13.640 800.000 14.240 ;
    END
  END sram_addr_b[6]
  PIN sram_addr_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END sram_addr_b[7]
  PIN sram_csb_a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END sram_csb_a
  PIN sram_csb_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END sram_csb_b
  PIN sram_din_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END sram_din_b[0]
  PIN sram_din_b[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1128.840 800.000 1129.440 ;
    END
  END sram_din_b[10]
  PIN sram_din_b[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END sram_din_b[11]
  PIN sram_din_b[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END sram_din_b[12]
  PIN sram_din_b[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1397.440 800.000 1398.040 ;
    END
  END sram_din_b[13]
  PIN sram_din_b[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 1596.000 116.290 1600.000 ;
    END
  END sram_din_b[14]
  PIN sram_din_b[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END sram_din_b[15]
  PIN sram_din_b[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END sram_din_b[16]
  PIN sram_din_b[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END sram_din_b[17]
  PIN sram_din_b[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 717.440 800.000 718.040 ;
    END
  END sram_din_b[18]
  PIN sram_din_b[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END sram_din_b[19]
  PIN sram_din_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END sram_din_b[1]
  PIN sram_din_b[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 683.440 800.000 684.040 ;
    END
  END sram_din_b[20]
  PIN sram_din_b[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 1596.000 705.550 1600.000 ;
    END
  END sram_din_b[21]
  PIN sram_din_b[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1033.640 800.000 1034.240 ;
    END
  END sram_din_b[22]
  PIN sram_din_b[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END sram_din_b[23]
  PIN sram_din_b[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 931.640 800.000 932.240 ;
    END
  END sram_din_b[24]
  PIN sram_din_b[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 74.840 800.000 75.440 ;
    END
  END sram_din_b[25]
  PIN sram_din_b[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1596.000 473.710 1600.000 ;
    END
  END sram_din_b[26]
  PIN sram_din_b[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END sram_din_b[27]
  PIN sram_din_b[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1193.440 800.000 1194.040 ;
    END
  END sram_din_b[28]
  PIN sram_din_b[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 1596.000 628.270 1600.000 ;
    END
  END sram_din_b[29]
  PIN sram_din_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 1596.000 486.590 1600.000 ;
    END
  END sram_din_b[2]
  PIN sram_din_b[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END sram_din_b[30]
  PIN sram_din_b[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 1596.000 641.150 1600.000 ;
    END
  END sram_din_b[31]
  PIN sram_din_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END sram_din_b[3]
  PIN sram_din_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END sram_din_b[4]
  PIN sram_din_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 561.040 800.000 561.640 ;
    END
  END sram_din_b[5]
  PIN sram_din_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 890.840 800.000 891.440 ;
    END
  END sram_din_b[6]
  PIN sram_din_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1227.440 800.000 1228.040 ;
    END
  END sram_din_b[7]
  PIN sram_din_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1596.000 10.030 1600.000 ;
    END
  END sram_din_b[8]
  PIN sram_din_b[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 170.040 800.000 170.640 ;
    END
  END sram_din_b[9]
  PIN sram_dout_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END sram_dout_a[0]
  PIN sram_dout_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1349.840 800.000 1350.440 ;
    END
  END sram_dout_a[10]
  PIN sram_dout_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END sram_dout_a[11]
  PIN sram_dout_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END sram_dout_a[12]
  PIN sram_dout_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 367.240 800.000 367.840 ;
    END
  END sram_dout_a[13]
  PIN sram_dout_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1596.000 744.190 1600.000 ;
    END
  END sram_dout_a[14]
  PIN sram_dout_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 319.640 800.000 320.240 ;
    END
  END sram_dout_a[15]
  PIN sram_dout_a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 547.440 800.000 548.040 ;
    END
  END sram_dout_a[16]
  PIN sram_dout_a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END sram_dout_a[17]
  PIN sram_dout_a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END sram_dout_a[18]
  PIN sram_dout_a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 397.840 800.000 398.440 ;
    END
  END sram_dout_a[19]
  PIN sram_dout_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 856.840 800.000 857.440 ;
    END
  END sram_dout_a[1]
  PIN sram_dout_a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1519.840 800.000 1520.440 ;
    END
  END sram_dout_a[20]
  PIN sram_dout_a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1596.000 51.890 1600.000 ;
    END
  END sram_dout_a[21]
  PIN sram_dout_a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 1596.000 3.590 1600.000 ;
    END
  END sram_dout_a[22]
  PIN sram_dout_a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.840 4.000 1401.440 ;
    END
  END sram_dout_a[23]
  PIN sram_dout_a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END sram_dout_a[24]
  PIN sram_dout_a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END sram_dout_a[25]
  PIN sram_dout_a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 527.040 800.000 527.640 ;
    END
  END sram_dout_a[26]
  PIN sram_dout_a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END sram_dout_a[27]
  PIN sram_dout_a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END sram_dout_a[28]
  PIN sram_dout_a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1492.640 800.000 1493.240 ;
    END
  END sram_dout_a[29]
  PIN sram_dout_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END sram_dout_a[2]
  PIN sram_dout_a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1596.000 219.330 1600.000 ;
    END
  END sram_dout_a[30]
  PIN sram_dout_a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END sram_dout_a[31]
  PIN sram_dout_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1596.000 499.470 1600.000 ;
    END
  END sram_dout_a[3]
  PIN sram_dout_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 1596.000 512.350 1600.000 ;
    END
  END sram_dout_a[4]
  PIN sram_dout_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END sram_dout_a[5]
  PIN sram_dout_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1596.000 103.410 1600.000 ;
    END
  END sram_dout_a[6]
  PIN sram_dout_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END sram_dout_a[7]
  PIN sram_dout_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END sram_dout_a[8]
  PIN sram_dout_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 306.040 800.000 306.640 ;
    END
  END sram_dout_a[9]
  PIN sram_dout_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END sram_dout_b[0]
  PIN sram_dout_b[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 710.640 800.000 711.240 ;
    END
  END sram_dout_b[10]
  PIN sram_dout_b[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END sram_dout_b[11]
  PIN sram_dout_b[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 822.840 800.000 823.440 ;
    END
  END sram_dout_b[12]
  PIN sram_dout_b[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END sram_dout_b[13]
  PIN sram_dout_b[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END sram_dout_b[14]
  PIN sram_dout_b[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END sram_dout_b[15]
  PIN sram_dout_b[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END sram_dout_b[16]
  PIN sram_dout_b[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1596.000 90.530 1600.000 ;
    END
  END sram_dout_b[17]
  PIN sram_dout_b[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 333.240 800.000 333.840 ;
    END
  END sram_dout_b[18]
  PIN sram_dout_b[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END sram_dout_b[19]
  PIN sram_dout_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 258.440 800.000 259.040 ;
    END
  END sram_dout_b[1]
  PIN sram_dout_b[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1329.440 800.000 1330.040 ;
    END
  END sram_dout_b[20]
  PIN sram_dout_b[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1594.640 800.000 1595.240 ;
    END
  END sram_dout_b[21]
  PIN sram_dout_b[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 278.840 800.000 279.440 ;
    END
  END sram_dout_b[22]
  PIN sram_dout_b[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END sram_dout_b[23]
  PIN sram_dout_b[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 595.040 800.000 595.640 ;
    END
  END sram_dout_b[24]
  PIN sram_dout_b[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1526.640 800.000 1527.240 ;
    END
  END sram_dout_b[25]
  PIN sram_dout_b[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END sram_dout_b[26]
  PIN sram_dout_b[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1343.040 800.000 1343.640 ;
    END
  END sram_dout_b[27]
  PIN sram_dout_b[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 251.640 800.000 252.240 ;
    END
  END sram_dout_b[28]
  PIN sram_dout_b[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END sram_dout_b[29]
  PIN sram_dout_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 737.840 800.000 738.440 ;
    END
  END sram_dout_b[2]
  PIN sram_dout_b[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1441.640 4.000 1442.240 ;
    END
  END sram_dout_b[30]
  PIN sram_dout_b[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END sram_dout_b[31]
  PIN sram_dout_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END sram_dout_b[3]
  PIN sram_dout_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END sram_dout_b[4]
  PIN sram_dout_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END sram_dout_b[5]
  PIN sram_dout_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END sram_dout_b[6]
  PIN sram_dout_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1506.240 800.000 1506.840 ;
    END
  END sram_dout_b[7]
  PIN sram_dout_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END sram_dout_b[8]
  PIN sram_dout_b[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END sram_dout_b[9]
  PIN sram_mask_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END sram_mask_b[0]
  PIN sram_mask_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 1596.000 257.970 1600.000 ;
    END
  END sram_mask_b[1]
  PIN sram_mask_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1596.000 763.510 1600.000 ;
    END
  END sram_mask_b[2]
  PIN sram_mask_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END sram_mask_b[3]
  PIN sram_web_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END sram_web_b
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 794.420 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 794.420 181.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 794.420 334.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 794.420 487.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 794.420 640.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 792.390 794.420 793.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 945.570 794.420 947.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1098.750 794.420 1100.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1251.930 794.420 1253.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1405.110 794.420 1406.710 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1558.290 794.420 1559.890 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1588.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 794.420 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 794.420 257.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 794.420 411.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 794.420 564.220 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 715.800 794.420 717.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 868.980 794.420 870.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1022.160 794.420 1023.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1175.340 794.420 1176.940 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1328.520 794.420 1330.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1481.700 794.420 1483.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1588.720 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 802.440 800.000 803.040 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1040.440 800.000 1041.040 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1596.000 32.570 1600.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1560.640 800.000 1561.240 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1472.240 800.000 1472.840 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 34.040 800.000 34.640 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1363.440 800.000 1364.040 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 965.640 800.000 966.240 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 479.440 800.000 480.040 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1596.000 58.330 1600.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1596.000 428.630 1600.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 265.240 800.000 265.840 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 4.000 1285.840 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1295.440 800.000 1296.040 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 1596.000 608.950 1600.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 1596.000 296.610 1600.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1074.440 800.000 1075.040 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 204.040 800.000 204.640 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1596.000 283.730 1600.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 163.240 800.000 163.840 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 850.040 800.000 850.640 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1596.000 757.070 1600.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 1596.000 232.210 1600.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 1596.000 538.110 1600.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1254.640 800.000 1255.240 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 1596.000 589.630 1600.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1479.040 800.000 1479.640 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 884.040 800.000 884.640 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 54.440 800.000 55.040 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1596.000 454.390 1600.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1234.240 800.000 1234.840 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 217.640 800.000 218.240 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 829.640 800.000 830.240 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 493.040 800.000 493.640 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 992.840 800.000 993.440 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1596.000 441.510 1600.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1581.040 800.000 1581.640 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 499.840 800.000 500.440 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1162.840 800.000 1163.440 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1596.000 798.930 1600.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1596.000 415.750 1600.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 574.640 800.000 575.240 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 6.840 800.000 7.440 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 0.040 800.000 0.640 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 149.640 800.000 150.240 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1596.000 180.690 1600.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1596.000 399.650 1600.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 751.440 800.000 752.040 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1356.640 800.000 1357.240 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1302.240 800.000 1302.840 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1596.000 380.330 1600.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1596.000 367.450 1600.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 40.840 800.000 41.440 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 979.240 800.000 979.840 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 1588.565 ;
      LAYER met1 ;
        RECT 0.070 10.640 798.950 1588.720 ;
      LAYER met2 ;
        RECT 0.100 1595.720 3.030 1598.525 ;
        RECT 3.870 1595.720 9.470 1598.525 ;
        RECT 10.310 1595.720 15.910 1598.525 ;
        RECT 16.750 1595.720 22.350 1598.525 ;
        RECT 23.190 1595.720 25.570 1598.525 ;
        RECT 26.410 1595.720 32.010 1598.525 ;
        RECT 32.850 1595.720 38.450 1598.525 ;
        RECT 39.290 1595.720 44.890 1598.525 ;
        RECT 45.730 1595.720 51.330 1598.525 ;
        RECT 52.170 1595.720 57.770 1598.525 ;
        RECT 58.610 1595.720 64.210 1598.525 ;
        RECT 65.050 1595.720 70.650 1598.525 ;
        RECT 71.490 1595.720 77.090 1598.525 ;
        RECT 77.930 1595.720 83.530 1598.525 ;
        RECT 84.370 1595.720 89.970 1598.525 ;
        RECT 90.810 1595.720 96.410 1598.525 ;
        RECT 97.250 1595.720 102.850 1598.525 ;
        RECT 103.690 1595.720 109.290 1598.525 ;
        RECT 110.130 1595.720 115.730 1598.525 ;
        RECT 116.570 1595.720 122.170 1598.525 ;
        RECT 123.010 1595.720 128.610 1598.525 ;
        RECT 129.450 1595.720 135.050 1598.525 ;
        RECT 135.890 1595.720 141.490 1598.525 ;
        RECT 142.330 1595.720 147.930 1598.525 ;
        RECT 148.770 1595.720 154.370 1598.525 ;
        RECT 155.210 1595.720 160.810 1598.525 ;
        RECT 161.650 1595.720 167.250 1598.525 ;
        RECT 168.090 1595.720 173.690 1598.525 ;
        RECT 174.530 1595.720 180.130 1598.525 ;
        RECT 180.970 1595.720 186.570 1598.525 ;
        RECT 187.410 1595.720 193.010 1598.525 ;
        RECT 193.850 1595.720 199.450 1598.525 ;
        RECT 200.290 1595.720 205.890 1598.525 ;
        RECT 206.730 1595.720 212.330 1598.525 ;
        RECT 213.170 1595.720 218.770 1598.525 ;
        RECT 219.610 1595.720 225.210 1598.525 ;
        RECT 226.050 1595.720 231.650 1598.525 ;
        RECT 232.490 1595.720 238.090 1598.525 ;
        RECT 238.930 1595.720 244.530 1598.525 ;
        RECT 245.370 1595.720 250.970 1598.525 ;
        RECT 251.810 1595.720 257.410 1598.525 ;
        RECT 258.250 1595.720 263.850 1598.525 ;
        RECT 264.690 1595.720 270.290 1598.525 ;
        RECT 271.130 1595.720 276.730 1598.525 ;
        RECT 277.570 1595.720 283.170 1598.525 ;
        RECT 284.010 1595.720 289.610 1598.525 ;
        RECT 290.450 1595.720 296.050 1598.525 ;
        RECT 296.890 1595.720 302.490 1598.525 ;
        RECT 303.330 1595.720 308.930 1598.525 ;
        RECT 309.770 1595.720 315.370 1598.525 ;
        RECT 316.210 1595.720 321.810 1598.525 ;
        RECT 322.650 1595.720 328.250 1598.525 ;
        RECT 329.090 1595.720 334.690 1598.525 ;
        RECT 335.530 1595.720 341.130 1598.525 ;
        RECT 341.970 1595.720 347.570 1598.525 ;
        RECT 348.410 1595.720 354.010 1598.525 ;
        RECT 354.850 1595.720 360.450 1598.525 ;
        RECT 361.290 1595.720 366.890 1598.525 ;
        RECT 367.730 1595.720 373.330 1598.525 ;
        RECT 374.170 1595.720 379.770 1598.525 ;
        RECT 380.610 1595.720 386.210 1598.525 ;
        RECT 387.050 1595.720 392.650 1598.525 ;
        RECT 393.490 1595.720 399.090 1598.525 ;
        RECT 399.930 1595.720 405.530 1598.525 ;
        RECT 406.370 1595.720 411.970 1598.525 ;
        RECT 412.810 1595.720 415.190 1598.525 ;
        RECT 416.030 1595.720 421.630 1598.525 ;
        RECT 422.470 1595.720 428.070 1598.525 ;
        RECT 428.910 1595.720 434.510 1598.525 ;
        RECT 435.350 1595.720 440.950 1598.525 ;
        RECT 441.790 1595.720 447.390 1598.525 ;
        RECT 448.230 1595.720 453.830 1598.525 ;
        RECT 454.670 1595.720 460.270 1598.525 ;
        RECT 461.110 1595.720 466.710 1598.525 ;
        RECT 467.550 1595.720 473.150 1598.525 ;
        RECT 473.990 1595.720 479.590 1598.525 ;
        RECT 480.430 1595.720 486.030 1598.525 ;
        RECT 486.870 1595.720 492.470 1598.525 ;
        RECT 493.310 1595.720 498.910 1598.525 ;
        RECT 499.750 1595.720 505.350 1598.525 ;
        RECT 506.190 1595.720 511.790 1598.525 ;
        RECT 512.630 1595.720 518.230 1598.525 ;
        RECT 519.070 1595.720 524.670 1598.525 ;
        RECT 525.510 1595.720 531.110 1598.525 ;
        RECT 531.950 1595.720 537.550 1598.525 ;
        RECT 538.390 1595.720 543.990 1598.525 ;
        RECT 544.830 1595.720 550.430 1598.525 ;
        RECT 551.270 1595.720 556.870 1598.525 ;
        RECT 557.710 1595.720 563.310 1598.525 ;
        RECT 564.150 1595.720 569.750 1598.525 ;
        RECT 570.590 1595.720 576.190 1598.525 ;
        RECT 577.030 1595.720 582.630 1598.525 ;
        RECT 583.470 1595.720 589.070 1598.525 ;
        RECT 589.910 1595.720 595.510 1598.525 ;
        RECT 596.350 1595.720 601.950 1598.525 ;
        RECT 602.790 1595.720 608.390 1598.525 ;
        RECT 609.230 1595.720 614.830 1598.525 ;
        RECT 615.670 1595.720 621.270 1598.525 ;
        RECT 622.110 1595.720 627.710 1598.525 ;
        RECT 628.550 1595.720 634.150 1598.525 ;
        RECT 634.990 1595.720 640.590 1598.525 ;
        RECT 641.430 1595.720 647.030 1598.525 ;
        RECT 647.870 1595.720 653.470 1598.525 ;
        RECT 654.310 1595.720 659.910 1598.525 ;
        RECT 660.750 1595.720 666.350 1598.525 ;
        RECT 667.190 1595.720 672.790 1598.525 ;
        RECT 673.630 1595.720 679.230 1598.525 ;
        RECT 680.070 1595.720 685.670 1598.525 ;
        RECT 686.510 1595.720 692.110 1598.525 ;
        RECT 692.950 1595.720 698.550 1598.525 ;
        RECT 699.390 1595.720 704.990 1598.525 ;
        RECT 705.830 1595.720 711.430 1598.525 ;
        RECT 712.270 1595.720 717.870 1598.525 ;
        RECT 718.710 1595.720 724.310 1598.525 ;
        RECT 725.150 1595.720 730.750 1598.525 ;
        RECT 731.590 1595.720 737.190 1598.525 ;
        RECT 738.030 1595.720 743.630 1598.525 ;
        RECT 744.470 1595.720 750.070 1598.525 ;
        RECT 750.910 1595.720 756.510 1598.525 ;
        RECT 757.350 1595.720 762.950 1598.525 ;
        RECT 763.790 1595.720 769.390 1598.525 ;
        RECT 770.230 1595.720 775.830 1598.525 ;
        RECT 776.670 1595.720 782.270 1598.525 ;
        RECT 783.110 1595.720 788.710 1598.525 ;
        RECT 789.550 1595.720 795.150 1598.525 ;
        RECT 795.990 1595.720 798.370 1598.525 ;
        RECT 0.100 4.280 798.920 1595.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 9.470 4.280 ;
        RECT 10.310 0.155 15.910 4.280 ;
        RECT 16.750 0.155 22.350 4.280 ;
        RECT 23.190 0.155 28.790 4.280 ;
        RECT 29.630 0.155 35.230 4.280 ;
        RECT 36.070 0.155 41.670 4.280 ;
        RECT 42.510 0.155 48.110 4.280 ;
        RECT 48.950 0.155 54.550 4.280 ;
        RECT 55.390 0.155 60.990 4.280 ;
        RECT 61.830 0.155 67.430 4.280 ;
        RECT 68.270 0.155 73.870 4.280 ;
        RECT 74.710 0.155 80.310 4.280 ;
        RECT 81.150 0.155 86.750 4.280 ;
        RECT 87.590 0.155 93.190 4.280 ;
        RECT 94.030 0.155 99.630 4.280 ;
        RECT 100.470 0.155 106.070 4.280 ;
        RECT 106.910 0.155 112.510 4.280 ;
        RECT 113.350 0.155 118.950 4.280 ;
        RECT 119.790 0.155 125.390 4.280 ;
        RECT 126.230 0.155 131.830 4.280 ;
        RECT 132.670 0.155 138.270 4.280 ;
        RECT 139.110 0.155 144.710 4.280 ;
        RECT 145.550 0.155 151.150 4.280 ;
        RECT 151.990 0.155 157.590 4.280 ;
        RECT 158.430 0.155 164.030 4.280 ;
        RECT 164.870 0.155 170.470 4.280 ;
        RECT 171.310 0.155 176.910 4.280 ;
        RECT 177.750 0.155 183.350 4.280 ;
        RECT 184.190 0.155 189.790 4.280 ;
        RECT 190.630 0.155 196.230 4.280 ;
        RECT 197.070 0.155 202.670 4.280 ;
        RECT 203.510 0.155 209.110 4.280 ;
        RECT 209.950 0.155 215.550 4.280 ;
        RECT 216.390 0.155 221.990 4.280 ;
        RECT 222.830 0.155 228.430 4.280 ;
        RECT 229.270 0.155 234.870 4.280 ;
        RECT 235.710 0.155 241.310 4.280 ;
        RECT 242.150 0.155 247.750 4.280 ;
        RECT 248.590 0.155 254.190 4.280 ;
        RECT 255.030 0.155 260.630 4.280 ;
        RECT 261.470 0.155 267.070 4.280 ;
        RECT 267.910 0.155 273.510 4.280 ;
        RECT 274.350 0.155 279.950 4.280 ;
        RECT 280.790 0.155 286.390 4.280 ;
        RECT 287.230 0.155 292.830 4.280 ;
        RECT 293.670 0.155 299.270 4.280 ;
        RECT 300.110 0.155 305.710 4.280 ;
        RECT 306.550 0.155 312.150 4.280 ;
        RECT 312.990 0.155 318.590 4.280 ;
        RECT 319.430 0.155 325.030 4.280 ;
        RECT 325.870 0.155 331.470 4.280 ;
        RECT 332.310 0.155 337.910 4.280 ;
        RECT 338.750 0.155 344.350 4.280 ;
        RECT 345.190 0.155 350.790 4.280 ;
        RECT 351.630 0.155 357.230 4.280 ;
        RECT 358.070 0.155 363.670 4.280 ;
        RECT 364.510 0.155 370.110 4.280 ;
        RECT 370.950 0.155 376.550 4.280 ;
        RECT 377.390 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 392.650 4.280 ;
        RECT 393.490 0.155 399.090 4.280 ;
        RECT 399.930 0.155 405.530 4.280 ;
        RECT 406.370 0.155 411.970 4.280 ;
        RECT 412.810 0.155 418.410 4.280 ;
        RECT 419.250 0.155 424.850 4.280 ;
        RECT 425.690 0.155 431.290 4.280 ;
        RECT 432.130 0.155 437.730 4.280 ;
        RECT 438.570 0.155 444.170 4.280 ;
        RECT 445.010 0.155 450.610 4.280 ;
        RECT 451.450 0.155 457.050 4.280 ;
        RECT 457.890 0.155 463.490 4.280 ;
        RECT 464.330 0.155 469.930 4.280 ;
        RECT 470.770 0.155 476.370 4.280 ;
        RECT 477.210 0.155 482.810 4.280 ;
        RECT 483.650 0.155 489.250 4.280 ;
        RECT 490.090 0.155 495.690 4.280 ;
        RECT 496.530 0.155 502.130 4.280 ;
        RECT 502.970 0.155 508.570 4.280 ;
        RECT 509.410 0.155 515.010 4.280 ;
        RECT 515.850 0.155 521.450 4.280 ;
        RECT 522.290 0.155 527.890 4.280 ;
        RECT 528.730 0.155 534.330 4.280 ;
        RECT 535.170 0.155 540.770 4.280 ;
        RECT 541.610 0.155 547.210 4.280 ;
        RECT 548.050 0.155 553.650 4.280 ;
        RECT 554.490 0.155 560.090 4.280 ;
        RECT 560.930 0.155 566.530 4.280 ;
        RECT 567.370 0.155 572.970 4.280 ;
        RECT 573.810 0.155 579.410 4.280 ;
        RECT 580.250 0.155 585.850 4.280 ;
        RECT 586.690 0.155 592.290 4.280 ;
        RECT 593.130 0.155 598.730 4.280 ;
        RECT 599.570 0.155 605.170 4.280 ;
        RECT 606.010 0.155 611.610 4.280 ;
        RECT 612.450 0.155 618.050 4.280 ;
        RECT 618.890 0.155 624.490 4.280 ;
        RECT 625.330 0.155 630.930 4.280 ;
        RECT 631.770 0.155 637.370 4.280 ;
        RECT 638.210 0.155 643.810 4.280 ;
        RECT 644.650 0.155 650.250 4.280 ;
        RECT 651.090 0.155 656.690 4.280 ;
        RECT 657.530 0.155 663.130 4.280 ;
        RECT 663.970 0.155 669.570 4.280 ;
        RECT 670.410 0.155 676.010 4.280 ;
        RECT 676.850 0.155 682.450 4.280 ;
        RECT 683.290 0.155 688.890 4.280 ;
        RECT 689.730 0.155 695.330 4.280 ;
        RECT 696.170 0.155 701.770 4.280 ;
        RECT 702.610 0.155 708.210 4.280 ;
        RECT 709.050 0.155 714.650 4.280 ;
        RECT 715.490 0.155 721.090 4.280 ;
        RECT 721.930 0.155 727.530 4.280 ;
        RECT 728.370 0.155 733.970 4.280 ;
        RECT 734.810 0.155 740.410 4.280 ;
        RECT 741.250 0.155 746.850 4.280 ;
        RECT 747.690 0.155 753.290 4.280 ;
        RECT 754.130 0.155 759.730 4.280 ;
        RECT 760.570 0.155 766.170 4.280 ;
        RECT 767.010 0.155 772.610 4.280 ;
        RECT 773.450 0.155 775.830 4.280 ;
        RECT 776.670 0.155 782.270 4.280 ;
        RECT 783.110 0.155 788.710 4.280 ;
        RECT 789.550 0.155 795.150 4.280 ;
        RECT 795.990 0.155 798.920 4.280 ;
      LAYER met3 ;
        RECT 4.400 1597.640 796.000 1598.505 ;
        RECT 4.000 1595.640 796.000 1597.640 ;
        RECT 4.000 1594.240 795.600 1595.640 ;
        RECT 4.000 1592.240 796.000 1594.240 ;
        RECT 4.400 1590.840 796.000 1592.240 ;
        RECT 4.000 1588.840 796.000 1590.840 ;
        RECT 4.000 1587.440 795.600 1588.840 ;
        RECT 4.000 1585.440 796.000 1587.440 ;
        RECT 4.400 1584.040 796.000 1585.440 ;
        RECT 4.000 1582.040 796.000 1584.040 ;
        RECT 4.000 1580.640 795.600 1582.040 ;
        RECT 4.000 1578.640 796.000 1580.640 ;
        RECT 4.400 1577.240 796.000 1578.640 ;
        RECT 4.000 1575.240 796.000 1577.240 ;
        RECT 4.000 1573.840 795.600 1575.240 ;
        RECT 4.000 1571.840 796.000 1573.840 ;
        RECT 4.400 1570.440 796.000 1571.840 ;
        RECT 4.000 1568.440 796.000 1570.440 ;
        RECT 4.000 1567.040 795.600 1568.440 ;
        RECT 4.000 1565.040 796.000 1567.040 ;
        RECT 4.400 1563.640 796.000 1565.040 ;
        RECT 4.000 1561.640 796.000 1563.640 ;
        RECT 4.000 1560.240 795.600 1561.640 ;
        RECT 4.000 1558.240 796.000 1560.240 ;
        RECT 4.400 1556.840 796.000 1558.240 ;
        RECT 4.000 1554.840 796.000 1556.840 ;
        RECT 4.000 1553.440 795.600 1554.840 ;
        RECT 4.000 1551.440 796.000 1553.440 ;
        RECT 4.400 1550.040 796.000 1551.440 ;
        RECT 4.000 1548.040 796.000 1550.040 ;
        RECT 4.000 1546.640 795.600 1548.040 ;
        RECT 4.000 1544.640 796.000 1546.640 ;
        RECT 4.400 1543.240 796.000 1544.640 ;
        RECT 4.000 1541.240 796.000 1543.240 ;
        RECT 4.000 1539.840 795.600 1541.240 ;
        RECT 4.000 1537.840 796.000 1539.840 ;
        RECT 4.400 1536.440 796.000 1537.840 ;
        RECT 4.000 1534.440 796.000 1536.440 ;
        RECT 4.000 1533.040 795.600 1534.440 ;
        RECT 4.000 1531.040 796.000 1533.040 ;
        RECT 4.400 1529.640 796.000 1531.040 ;
        RECT 4.000 1527.640 796.000 1529.640 ;
        RECT 4.000 1526.240 795.600 1527.640 ;
        RECT 4.000 1524.240 796.000 1526.240 ;
        RECT 4.400 1522.840 796.000 1524.240 ;
        RECT 4.000 1520.840 796.000 1522.840 ;
        RECT 4.000 1519.440 795.600 1520.840 ;
        RECT 4.000 1517.440 796.000 1519.440 ;
        RECT 4.400 1516.040 796.000 1517.440 ;
        RECT 4.000 1514.040 796.000 1516.040 ;
        RECT 4.000 1512.640 795.600 1514.040 ;
        RECT 4.000 1510.640 796.000 1512.640 ;
        RECT 4.400 1509.240 796.000 1510.640 ;
        RECT 4.000 1507.240 796.000 1509.240 ;
        RECT 4.000 1505.840 795.600 1507.240 ;
        RECT 4.000 1503.840 796.000 1505.840 ;
        RECT 4.400 1502.440 796.000 1503.840 ;
        RECT 4.000 1500.440 796.000 1502.440 ;
        RECT 4.000 1499.040 795.600 1500.440 ;
        RECT 4.000 1497.040 796.000 1499.040 ;
        RECT 4.400 1495.640 796.000 1497.040 ;
        RECT 4.000 1493.640 796.000 1495.640 ;
        RECT 4.000 1492.240 795.600 1493.640 ;
        RECT 4.000 1490.240 796.000 1492.240 ;
        RECT 4.400 1488.840 796.000 1490.240 ;
        RECT 4.000 1486.840 796.000 1488.840 ;
        RECT 4.000 1485.440 795.600 1486.840 ;
        RECT 4.000 1483.440 796.000 1485.440 ;
        RECT 4.400 1482.040 796.000 1483.440 ;
        RECT 4.000 1480.040 796.000 1482.040 ;
        RECT 4.000 1478.640 795.600 1480.040 ;
        RECT 4.000 1476.640 796.000 1478.640 ;
        RECT 4.400 1475.240 796.000 1476.640 ;
        RECT 4.000 1473.240 796.000 1475.240 ;
        RECT 4.000 1471.840 795.600 1473.240 ;
        RECT 4.000 1469.840 796.000 1471.840 ;
        RECT 4.400 1468.440 796.000 1469.840 ;
        RECT 4.000 1466.440 796.000 1468.440 ;
        RECT 4.000 1465.040 795.600 1466.440 ;
        RECT 4.000 1463.040 796.000 1465.040 ;
        RECT 4.400 1461.640 796.000 1463.040 ;
        RECT 4.000 1459.640 796.000 1461.640 ;
        RECT 4.000 1458.240 795.600 1459.640 ;
        RECT 4.000 1456.240 796.000 1458.240 ;
        RECT 4.400 1454.840 796.000 1456.240 ;
        RECT 4.000 1452.840 796.000 1454.840 ;
        RECT 4.000 1451.440 795.600 1452.840 ;
        RECT 4.000 1449.440 796.000 1451.440 ;
        RECT 4.400 1448.040 796.000 1449.440 ;
        RECT 4.000 1446.040 796.000 1448.040 ;
        RECT 4.000 1444.640 795.600 1446.040 ;
        RECT 4.000 1442.640 796.000 1444.640 ;
        RECT 4.400 1441.240 796.000 1442.640 ;
        RECT 4.000 1439.240 796.000 1441.240 ;
        RECT 4.000 1437.840 795.600 1439.240 ;
        RECT 4.000 1435.840 796.000 1437.840 ;
        RECT 4.400 1434.440 796.000 1435.840 ;
        RECT 4.000 1432.440 796.000 1434.440 ;
        RECT 4.000 1431.040 795.600 1432.440 ;
        RECT 4.000 1429.040 796.000 1431.040 ;
        RECT 4.400 1427.640 796.000 1429.040 ;
        RECT 4.000 1425.640 796.000 1427.640 ;
        RECT 4.000 1424.240 795.600 1425.640 ;
        RECT 4.000 1422.240 796.000 1424.240 ;
        RECT 4.400 1420.840 796.000 1422.240 ;
        RECT 4.000 1418.840 796.000 1420.840 ;
        RECT 4.000 1417.440 795.600 1418.840 ;
        RECT 4.000 1415.440 796.000 1417.440 ;
        RECT 4.400 1414.040 796.000 1415.440 ;
        RECT 4.000 1412.040 796.000 1414.040 ;
        RECT 4.000 1410.640 795.600 1412.040 ;
        RECT 4.000 1408.640 796.000 1410.640 ;
        RECT 4.400 1407.240 796.000 1408.640 ;
        RECT 4.000 1405.240 796.000 1407.240 ;
        RECT 4.000 1403.840 795.600 1405.240 ;
        RECT 4.000 1401.840 796.000 1403.840 ;
        RECT 4.400 1400.440 796.000 1401.840 ;
        RECT 4.000 1398.440 796.000 1400.440 ;
        RECT 4.000 1397.040 795.600 1398.440 ;
        RECT 4.000 1395.040 796.000 1397.040 ;
        RECT 4.400 1393.640 796.000 1395.040 ;
        RECT 4.000 1391.640 796.000 1393.640 ;
        RECT 4.000 1390.240 795.600 1391.640 ;
        RECT 4.000 1388.240 796.000 1390.240 ;
        RECT 4.400 1386.840 796.000 1388.240 ;
        RECT 4.000 1384.840 796.000 1386.840 ;
        RECT 4.000 1383.440 795.600 1384.840 ;
        RECT 4.000 1381.440 796.000 1383.440 ;
        RECT 4.400 1380.040 796.000 1381.440 ;
        RECT 4.000 1378.040 796.000 1380.040 ;
        RECT 4.000 1376.640 795.600 1378.040 ;
        RECT 4.000 1374.640 796.000 1376.640 ;
        RECT 4.400 1373.240 796.000 1374.640 ;
        RECT 4.000 1371.240 796.000 1373.240 ;
        RECT 4.000 1369.840 795.600 1371.240 ;
        RECT 4.000 1367.840 796.000 1369.840 ;
        RECT 4.400 1366.440 796.000 1367.840 ;
        RECT 4.000 1364.440 796.000 1366.440 ;
        RECT 4.000 1363.040 795.600 1364.440 ;
        RECT 4.000 1361.040 796.000 1363.040 ;
        RECT 4.400 1359.640 796.000 1361.040 ;
        RECT 4.000 1357.640 796.000 1359.640 ;
        RECT 4.000 1356.240 795.600 1357.640 ;
        RECT 4.000 1354.240 796.000 1356.240 ;
        RECT 4.400 1352.840 796.000 1354.240 ;
        RECT 4.000 1350.840 796.000 1352.840 ;
        RECT 4.000 1349.440 795.600 1350.840 ;
        RECT 4.000 1347.440 796.000 1349.440 ;
        RECT 4.400 1346.040 796.000 1347.440 ;
        RECT 4.000 1344.040 796.000 1346.040 ;
        RECT 4.000 1342.640 795.600 1344.040 ;
        RECT 4.000 1340.640 796.000 1342.640 ;
        RECT 4.400 1339.240 796.000 1340.640 ;
        RECT 4.000 1337.240 796.000 1339.240 ;
        RECT 4.000 1335.840 795.600 1337.240 ;
        RECT 4.000 1333.840 796.000 1335.840 ;
        RECT 4.400 1332.440 796.000 1333.840 ;
        RECT 4.000 1330.440 796.000 1332.440 ;
        RECT 4.000 1329.040 795.600 1330.440 ;
        RECT 4.000 1327.040 796.000 1329.040 ;
        RECT 4.400 1325.640 796.000 1327.040 ;
        RECT 4.000 1323.640 796.000 1325.640 ;
        RECT 4.000 1322.240 795.600 1323.640 ;
        RECT 4.000 1320.240 796.000 1322.240 ;
        RECT 4.400 1318.840 796.000 1320.240 ;
        RECT 4.000 1316.840 796.000 1318.840 ;
        RECT 4.000 1315.440 795.600 1316.840 ;
        RECT 4.000 1313.440 796.000 1315.440 ;
        RECT 4.400 1312.040 796.000 1313.440 ;
        RECT 4.000 1310.040 796.000 1312.040 ;
        RECT 4.000 1308.640 795.600 1310.040 ;
        RECT 4.000 1306.640 796.000 1308.640 ;
        RECT 4.400 1305.240 796.000 1306.640 ;
        RECT 4.000 1303.240 796.000 1305.240 ;
        RECT 4.000 1301.840 795.600 1303.240 ;
        RECT 4.000 1299.840 796.000 1301.840 ;
        RECT 4.400 1298.440 796.000 1299.840 ;
        RECT 4.000 1296.440 796.000 1298.440 ;
        RECT 4.000 1295.040 795.600 1296.440 ;
        RECT 4.000 1293.040 796.000 1295.040 ;
        RECT 4.400 1291.640 796.000 1293.040 ;
        RECT 4.000 1289.640 796.000 1291.640 ;
        RECT 4.000 1288.240 795.600 1289.640 ;
        RECT 4.000 1286.240 796.000 1288.240 ;
        RECT 4.400 1284.840 796.000 1286.240 ;
        RECT 4.000 1282.840 796.000 1284.840 ;
        RECT 4.000 1281.440 795.600 1282.840 ;
        RECT 4.000 1279.440 796.000 1281.440 ;
        RECT 4.400 1278.040 796.000 1279.440 ;
        RECT 4.000 1276.040 796.000 1278.040 ;
        RECT 4.000 1274.640 795.600 1276.040 ;
        RECT 4.000 1272.640 796.000 1274.640 ;
        RECT 4.400 1271.240 796.000 1272.640 ;
        RECT 4.000 1269.240 796.000 1271.240 ;
        RECT 4.000 1267.840 795.600 1269.240 ;
        RECT 4.000 1265.840 796.000 1267.840 ;
        RECT 4.400 1264.440 796.000 1265.840 ;
        RECT 4.000 1262.440 796.000 1264.440 ;
        RECT 4.000 1261.040 795.600 1262.440 ;
        RECT 4.000 1259.040 796.000 1261.040 ;
        RECT 4.400 1257.640 796.000 1259.040 ;
        RECT 4.000 1255.640 796.000 1257.640 ;
        RECT 4.000 1254.240 795.600 1255.640 ;
        RECT 4.000 1252.240 796.000 1254.240 ;
        RECT 4.400 1250.840 796.000 1252.240 ;
        RECT 4.000 1248.840 796.000 1250.840 ;
        RECT 4.000 1247.440 795.600 1248.840 ;
        RECT 4.000 1245.440 796.000 1247.440 ;
        RECT 4.400 1244.040 796.000 1245.440 ;
        RECT 4.000 1242.040 796.000 1244.040 ;
        RECT 4.000 1240.640 795.600 1242.040 ;
        RECT 4.000 1238.640 796.000 1240.640 ;
        RECT 4.400 1237.240 796.000 1238.640 ;
        RECT 4.000 1235.240 796.000 1237.240 ;
        RECT 4.000 1233.840 795.600 1235.240 ;
        RECT 4.000 1231.840 796.000 1233.840 ;
        RECT 4.400 1230.440 796.000 1231.840 ;
        RECT 4.000 1228.440 796.000 1230.440 ;
        RECT 4.000 1227.040 795.600 1228.440 ;
        RECT 4.000 1225.040 796.000 1227.040 ;
        RECT 4.400 1223.640 796.000 1225.040 ;
        RECT 4.000 1221.640 796.000 1223.640 ;
        RECT 4.400 1220.240 795.600 1221.640 ;
        RECT 4.000 1214.840 796.000 1220.240 ;
        RECT 4.400 1213.440 795.600 1214.840 ;
        RECT 4.000 1208.040 796.000 1213.440 ;
        RECT 4.400 1206.640 795.600 1208.040 ;
        RECT 4.000 1201.240 796.000 1206.640 ;
        RECT 4.400 1199.840 795.600 1201.240 ;
        RECT 4.000 1194.440 796.000 1199.840 ;
        RECT 4.400 1193.040 795.600 1194.440 ;
        RECT 4.000 1191.040 796.000 1193.040 ;
        RECT 4.000 1189.640 795.600 1191.040 ;
        RECT 4.000 1187.640 796.000 1189.640 ;
        RECT 4.400 1186.240 796.000 1187.640 ;
        RECT 4.000 1184.240 796.000 1186.240 ;
        RECT 4.000 1182.840 795.600 1184.240 ;
        RECT 4.000 1180.840 796.000 1182.840 ;
        RECT 4.400 1179.440 796.000 1180.840 ;
        RECT 4.000 1177.440 796.000 1179.440 ;
        RECT 4.000 1176.040 795.600 1177.440 ;
        RECT 4.000 1174.040 796.000 1176.040 ;
        RECT 4.400 1172.640 796.000 1174.040 ;
        RECT 4.000 1170.640 796.000 1172.640 ;
        RECT 4.000 1169.240 795.600 1170.640 ;
        RECT 4.000 1167.240 796.000 1169.240 ;
        RECT 4.400 1165.840 796.000 1167.240 ;
        RECT 4.000 1163.840 796.000 1165.840 ;
        RECT 4.000 1162.440 795.600 1163.840 ;
        RECT 4.000 1160.440 796.000 1162.440 ;
        RECT 4.400 1159.040 796.000 1160.440 ;
        RECT 4.000 1157.040 796.000 1159.040 ;
        RECT 4.000 1155.640 795.600 1157.040 ;
        RECT 4.000 1153.640 796.000 1155.640 ;
        RECT 4.400 1152.240 796.000 1153.640 ;
        RECT 4.000 1150.240 796.000 1152.240 ;
        RECT 4.000 1148.840 795.600 1150.240 ;
        RECT 4.000 1146.840 796.000 1148.840 ;
        RECT 4.400 1145.440 796.000 1146.840 ;
        RECT 4.000 1143.440 796.000 1145.440 ;
        RECT 4.000 1142.040 795.600 1143.440 ;
        RECT 4.000 1140.040 796.000 1142.040 ;
        RECT 4.400 1138.640 796.000 1140.040 ;
        RECT 4.000 1136.640 796.000 1138.640 ;
        RECT 4.000 1135.240 795.600 1136.640 ;
        RECT 4.000 1133.240 796.000 1135.240 ;
        RECT 4.400 1131.840 796.000 1133.240 ;
        RECT 4.000 1129.840 796.000 1131.840 ;
        RECT 4.000 1128.440 795.600 1129.840 ;
        RECT 4.000 1126.440 796.000 1128.440 ;
        RECT 4.400 1125.040 796.000 1126.440 ;
        RECT 4.000 1123.040 796.000 1125.040 ;
        RECT 4.000 1121.640 795.600 1123.040 ;
        RECT 4.000 1119.640 796.000 1121.640 ;
        RECT 4.400 1118.240 796.000 1119.640 ;
        RECT 4.000 1116.240 796.000 1118.240 ;
        RECT 4.000 1114.840 795.600 1116.240 ;
        RECT 4.000 1112.840 796.000 1114.840 ;
        RECT 4.400 1111.440 796.000 1112.840 ;
        RECT 4.000 1109.440 796.000 1111.440 ;
        RECT 4.000 1108.040 795.600 1109.440 ;
        RECT 4.000 1106.040 796.000 1108.040 ;
        RECT 4.400 1104.640 796.000 1106.040 ;
        RECT 4.000 1102.640 796.000 1104.640 ;
        RECT 4.000 1101.240 795.600 1102.640 ;
        RECT 4.000 1099.240 796.000 1101.240 ;
        RECT 4.400 1097.840 796.000 1099.240 ;
        RECT 4.000 1095.840 796.000 1097.840 ;
        RECT 4.000 1094.440 795.600 1095.840 ;
        RECT 4.000 1092.440 796.000 1094.440 ;
        RECT 4.400 1091.040 796.000 1092.440 ;
        RECT 4.000 1089.040 796.000 1091.040 ;
        RECT 4.000 1087.640 795.600 1089.040 ;
        RECT 4.000 1085.640 796.000 1087.640 ;
        RECT 4.400 1084.240 796.000 1085.640 ;
        RECT 4.000 1082.240 796.000 1084.240 ;
        RECT 4.000 1080.840 795.600 1082.240 ;
        RECT 4.000 1078.840 796.000 1080.840 ;
        RECT 4.400 1077.440 796.000 1078.840 ;
        RECT 4.000 1075.440 796.000 1077.440 ;
        RECT 4.000 1074.040 795.600 1075.440 ;
        RECT 4.000 1072.040 796.000 1074.040 ;
        RECT 4.400 1070.640 796.000 1072.040 ;
        RECT 4.000 1068.640 796.000 1070.640 ;
        RECT 4.000 1067.240 795.600 1068.640 ;
        RECT 4.000 1065.240 796.000 1067.240 ;
        RECT 4.400 1063.840 796.000 1065.240 ;
        RECT 4.000 1061.840 796.000 1063.840 ;
        RECT 4.000 1060.440 795.600 1061.840 ;
        RECT 4.000 1058.440 796.000 1060.440 ;
        RECT 4.400 1057.040 796.000 1058.440 ;
        RECT 4.000 1055.040 796.000 1057.040 ;
        RECT 4.000 1053.640 795.600 1055.040 ;
        RECT 4.000 1051.640 796.000 1053.640 ;
        RECT 4.400 1050.240 796.000 1051.640 ;
        RECT 4.000 1048.240 796.000 1050.240 ;
        RECT 4.000 1046.840 795.600 1048.240 ;
        RECT 4.000 1044.840 796.000 1046.840 ;
        RECT 4.400 1043.440 796.000 1044.840 ;
        RECT 4.000 1041.440 796.000 1043.440 ;
        RECT 4.000 1040.040 795.600 1041.440 ;
        RECT 4.000 1038.040 796.000 1040.040 ;
        RECT 4.400 1036.640 796.000 1038.040 ;
        RECT 4.000 1034.640 796.000 1036.640 ;
        RECT 4.000 1033.240 795.600 1034.640 ;
        RECT 4.000 1031.240 796.000 1033.240 ;
        RECT 4.400 1029.840 796.000 1031.240 ;
        RECT 4.000 1027.840 796.000 1029.840 ;
        RECT 4.000 1026.440 795.600 1027.840 ;
        RECT 4.000 1024.440 796.000 1026.440 ;
        RECT 4.400 1023.040 796.000 1024.440 ;
        RECT 4.000 1021.040 796.000 1023.040 ;
        RECT 4.000 1019.640 795.600 1021.040 ;
        RECT 4.000 1017.640 796.000 1019.640 ;
        RECT 4.400 1016.240 796.000 1017.640 ;
        RECT 4.000 1014.240 796.000 1016.240 ;
        RECT 4.000 1012.840 795.600 1014.240 ;
        RECT 4.000 1010.840 796.000 1012.840 ;
        RECT 4.400 1009.440 796.000 1010.840 ;
        RECT 4.000 1007.440 796.000 1009.440 ;
        RECT 4.000 1006.040 795.600 1007.440 ;
        RECT 4.000 1004.040 796.000 1006.040 ;
        RECT 4.400 1002.640 796.000 1004.040 ;
        RECT 4.000 1000.640 796.000 1002.640 ;
        RECT 4.000 999.240 795.600 1000.640 ;
        RECT 4.000 997.240 796.000 999.240 ;
        RECT 4.400 995.840 796.000 997.240 ;
        RECT 4.000 993.840 796.000 995.840 ;
        RECT 4.000 992.440 795.600 993.840 ;
        RECT 4.000 990.440 796.000 992.440 ;
        RECT 4.400 989.040 796.000 990.440 ;
        RECT 4.000 987.040 796.000 989.040 ;
        RECT 4.000 985.640 795.600 987.040 ;
        RECT 4.000 983.640 796.000 985.640 ;
        RECT 4.400 982.240 796.000 983.640 ;
        RECT 4.000 980.240 796.000 982.240 ;
        RECT 4.000 978.840 795.600 980.240 ;
        RECT 4.000 976.840 796.000 978.840 ;
        RECT 4.400 975.440 796.000 976.840 ;
        RECT 4.000 973.440 796.000 975.440 ;
        RECT 4.000 972.040 795.600 973.440 ;
        RECT 4.000 970.040 796.000 972.040 ;
        RECT 4.400 968.640 796.000 970.040 ;
        RECT 4.000 966.640 796.000 968.640 ;
        RECT 4.000 965.240 795.600 966.640 ;
        RECT 4.000 963.240 796.000 965.240 ;
        RECT 4.400 961.840 796.000 963.240 ;
        RECT 4.000 959.840 796.000 961.840 ;
        RECT 4.000 958.440 795.600 959.840 ;
        RECT 4.000 956.440 796.000 958.440 ;
        RECT 4.400 955.040 796.000 956.440 ;
        RECT 4.000 953.040 796.000 955.040 ;
        RECT 4.000 951.640 795.600 953.040 ;
        RECT 4.000 949.640 796.000 951.640 ;
        RECT 4.400 948.240 796.000 949.640 ;
        RECT 4.000 946.240 796.000 948.240 ;
        RECT 4.000 944.840 795.600 946.240 ;
        RECT 4.000 942.840 796.000 944.840 ;
        RECT 4.400 941.440 796.000 942.840 ;
        RECT 4.000 939.440 796.000 941.440 ;
        RECT 4.000 938.040 795.600 939.440 ;
        RECT 4.000 936.040 796.000 938.040 ;
        RECT 4.400 934.640 796.000 936.040 ;
        RECT 4.000 932.640 796.000 934.640 ;
        RECT 4.000 931.240 795.600 932.640 ;
        RECT 4.000 929.240 796.000 931.240 ;
        RECT 4.400 927.840 796.000 929.240 ;
        RECT 4.000 925.840 796.000 927.840 ;
        RECT 4.000 924.440 795.600 925.840 ;
        RECT 4.000 922.440 796.000 924.440 ;
        RECT 4.400 921.040 796.000 922.440 ;
        RECT 4.000 919.040 796.000 921.040 ;
        RECT 4.000 917.640 795.600 919.040 ;
        RECT 4.000 915.640 796.000 917.640 ;
        RECT 4.400 914.240 796.000 915.640 ;
        RECT 4.000 912.240 796.000 914.240 ;
        RECT 4.000 910.840 795.600 912.240 ;
        RECT 4.000 908.840 796.000 910.840 ;
        RECT 4.400 907.440 796.000 908.840 ;
        RECT 4.000 905.440 796.000 907.440 ;
        RECT 4.000 904.040 795.600 905.440 ;
        RECT 4.000 902.040 796.000 904.040 ;
        RECT 4.400 900.640 796.000 902.040 ;
        RECT 4.000 898.640 796.000 900.640 ;
        RECT 4.000 897.240 795.600 898.640 ;
        RECT 4.000 895.240 796.000 897.240 ;
        RECT 4.400 893.840 796.000 895.240 ;
        RECT 4.000 891.840 796.000 893.840 ;
        RECT 4.000 890.440 795.600 891.840 ;
        RECT 4.000 888.440 796.000 890.440 ;
        RECT 4.400 887.040 796.000 888.440 ;
        RECT 4.000 885.040 796.000 887.040 ;
        RECT 4.000 883.640 795.600 885.040 ;
        RECT 4.000 881.640 796.000 883.640 ;
        RECT 4.400 880.240 796.000 881.640 ;
        RECT 4.000 878.240 796.000 880.240 ;
        RECT 4.000 876.840 795.600 878.240 ;
        RECT 4.000 874.840 796.000 876.840 ;
        RECT 4.400 873.440 796.000 874.840 ;
        RECT 4.000 871.440 796.000 873.440 ;
        RECT 4.000 870.040 795.600 871.440 ;
        RECT 4.000 868.040 796.000 870.040 ;
        RECT 4.400 866.640 796.000 868.040 ;
        RECT 4.000 864.640 796.000 866.640 ;
        RECT 4.000 863.240 795.600 864.640 ;
        RECT 4.000 861.240 796.000 863.240 ;
        RECT 4.400 859.840 796.000 861.240 ;
        RECT 4.000 857.840 796.000 859.840 ;
        RECT 4.000 856.440 795.600 857.840 ;
        RECT 4.000 854.440 796.000 856.440 ;
        RECT 4.400 853.040 796.000 854.440 ;
        RECT 4.000 851.040 796.000 853.040 ;
        RECT 4.000 849.640 795.600 851.040 ;
        RECT 4.000 847.640 796.000 849.640 ;
        RECT 4.400 846.240 796.000 847.640 ;
        RECT 4.000 844.240 796.000 846.240 ;
        RECT 4.000 842.840 795.600 844.240 ;
        RECT 4.000 840.840 796.000 842.840 ;
        RECT 4.400 839.440 796.000 840.840 ;
        RECT 4.000 837.440 796.000 839.440 ;
        RECT 4.000 836.040 795.600 837.440 ;
        RECT 4.000 834.040 796.000 836.040 ;
        RECT 4.400 832.640 796.000 834.040 ;
        RECT 4.000 830.640 796.000 832.640 ;
        RECT 4.000 829.240 795.600 830.640 ;
        RECT 4.000 827.240 796.000 829.240 ;
        RECT 4.400 825.840 796.000 827.240 ;
        RECT 4.000 823.840 796.000 825.840 ;
        RECT 4.000 822.440 795.600 823.840 ;
        RECT 4.000 820.440 796.000 822.440 ;
        RECT 4.400 819.040 796.000 820.440 ;
        RECT 4.000 817.040 796.000 819.040 ;
        RECT 4.000 815.640 795.600 817.040 ;
        RECT 4.000 813.640 796.000 815.640 ;
        RECT 4.400 812.240 796.000 813.640 ;
        RECT 4.000 810.240 796.000 812.240 ;
        RECT 4.400 808.840 795.600 810.240 ;
        RECT 4.000 803.440 796.000 808.840 ;
        RECT 4.400 802.040 795.600 803.440 ;
        RECT 4.000 796.640 796.000 802.040 ;
        RECT 4.400 795.240 795.600 796.640 ;
        RECT 4.000 789.840 796.000 795.240 ;
        RECT 4.400 788.440 795.600 789.840 ;
        RECT 4.000 786.440 796.000 788.440 ;
        RECT 4.000 785.040 795.600 786.440 ;
        RECT 4.000 783.040 796.000 785.040 ;
        RECT 4.400 781.640 796.000 783.040 ;
        RECT 4.000 779.640 796.000 781.640 ;
        RECT 4.000 778.240 795.600 779.640 ;
        RECT 4.000 776.240 796.000 778.240 ;
        RECT 4.400 774.840 796.000 776.240 ;
        RECT 4.000 772.840 796.000 774.840 ;
        RECT 4.000 771.440 795.600 772.840 ;
        RECT 4.000 769.440 796.000 771.440 ;
        RECT 4.400 768.040 796.000 769.440 ;
        RECT 4.000 766.040 796.000 768.040 ;
        RECT 4.000 764.640 795.600 766.040 ;
        RECT 4.000 762.640 796.000 764.640 ;
        RECT 4.400 761.240 796.000 762.640 ;
        RECT 4.000 759.240 796.000 761.240 ;
        RECT 4.000 757.840 795.600 759.240 ;
        RECT 4.000 755.840 796.000 757.840 ;
        RECT 4.400 754.440 796.000 755.840 ;
        RECT 4.000 752.440 796.000 754.440 ;
        RECT 4.000 751.040 795.600 752.440 ;
        RECT 4.000 749.040 796.000 751.040 ;
        RECT 4.400 747.640 796.000 749.040 ;
        RECT 4.000 745.640 796.000 747.640 ;
        RECT 4.000 744.240 795.600 745.640 ;
        RECT 4.000 742.240 796.000 744.240 ;
        RECT 4.400 740.840 796.000 742.240 ;
        RECT 4.000 738.840 796.000 740.840 ;
        RECT 4.000 737.440 795.600 738.840 ;
        RECT 4.000 735.440 796.000 737.440 ;
        RECT 4.400 734.040 796.000 735.440 ;
        RECT 4.000 732.040 796.000 734.040 ;
        RECT 4.000 730.640 795.600 732.040 ;
        RECT 4.000 728.640 796.000 730.640 ;
        RECT 4.400 727.240 796.000 728.640 ;
        RECT 4.000 725.240 796.000 727.240 ;
        RECT 4.000 723.840 795.600 725.240 ;
        RECT 4.000 721.840 796.000 723.840 ;
        RECT 4.400 720.440 796.000 721.840 ;
        RECT 4.000 718.440 796.000 720.440 ;
        RECT 4.000 717.040 795.600 718.440 ;
        RECT 4.000 715.040 796.000 717.040 ;
        RECT 4.400 713.640 796.000 715.040 ;
        RECT 4.000 711.640 796.000 713.640 ;
        RECT 4.000 710.240 795.600 711.640 ;
        RECT 4.000 708.240 796.000 710.240 ;
        RECT 4.400 706.840 796.000 708.240 ;
        RECT 4.000 704.840 796.000 706.840 ;
        RECT 4.000 703.440 795.600 704.840 ;
        RECT 4.000 701.440 796.000 703.440 ;
        RECT 4.400 700.040 796.000 701.440 ;
        RECT 4.000 698.040 796.000 700.040 ;
        RECT 4.000 696.640 795.600 698.040 ;
        RECT 4.000 694.640 796.000 696.640 ;
        RECT 4.400 693.240 796.000 694.640 ;
        RECT 4.000 691.240 796.000 693.240 ;
        RECT 4.000 689.840 795.600 691.240 ;
        RECT 4.000 687.840 796.000 689.840 ;
        RECT 4.400 686.440 796.000 687.840 ;
        RECT 4.000 684.440 796.000 686.440 ;
        RECT 4.000 683.040 795.600 684.440 ;
        RECT 4.000 681.040 796.000 683.040 ;
        RECT 4.400 679.640 796.000 681.040 ;
        RECT 4.000 677.640 796.000 679.640 ;
        RECT 4.000 676.240 795.600 677.640 ;
        RECT 4.000 674.240 796.000 676.240 ;
        RECT 4.400 672.840 796.000 674.240 ;
        RECT 4.000 670.840 796.000 672.840 ;
        RECT 4.000 669.440 795.600 670.840 ;
        RECT 4.000 667.440 796.000 669.440 ;
        RECT 4.400 666.040 796.000 667.440 ;
        RECT 4.000 664.040 796.000 666.040 ;
        RECT 4.000 662.640 795.600 664.040 ;
        RECT 4.000 660.640 796.000 662.640 ;
        RECT 4.400 659.240 796.000 660.640 ;
        RECT 4.000 657.240 796.000 659.240 ;
        RECT 4.000 655.840 795.600 657.240 ;
        RECT 4.000 653.840 796.000 655.840 ;
        RECT 4.400 652.440 796.000 653.840 ;
        RECT 4.000 650.440 796.000 652.440 ;
        RECT 4.000 649.040 795.600 650.440 ;
        RECT 4.000 647.040 796.000 649.040 ;
        RECT 4.400 645.640 796.000 647.040 ;
        RECT 4.000 643.640 796.000 645.640 ;
        RECT 4.000 642.240 795.600 643.640 ;
        RECT 4.000 640.240 796.000 642.240 ;
        RECT 4.400 638.840 796.000 640.240 ;
        RECT 4.000 636.840 796.000 638.840 ;
        RECT 4.000 635.440 795.600 636.840 ;
        RECT 4.000 633.440 796.000 635.440 ;
        RECT 4.400 632.040 796.000 633.440 ;
        RECT 4.000 630.040 796.000 632.040 ;
        RECT 4.000 628.640 795.600 630.040 ;
        RECT 4.000 626.640 796.000 628.640 ;
        RECT 4.400 625.240 796.000 626.640 ;
        RECT 4.000 623.240 796.000 625.240 ;
        RECT 4.000 621.840 795.600 623.240 ;
        RECT 4.000 619.840 796.000 621.840 ;
        RECT 4.400 618.440 796.000 619.840 ;
        RECT 4.000 616.440 796.000 618.440 ;
        RECT 4.000 615.040 795.600 616.440 ;
        RECT 4.000 613.040 796.000 615.040 ;
        RECT 4.400 611.640 796.000 613.040 ;
        RECT 4.000 609.640 796.000 611.640 ;
        RECT 4.000 608.240 795.600 609.640 ;
        RECT 4.000 606.240 796.000 608.240 ;
        RECT 4.400 604.840 796.000 606.240 ;
        RECT 4.000 602.840 796.000 604.840 ;
        RECT 4.000 601.440 795.600 602.840 ;
        RECT 4.000 599.440 796.000 601.440 ;
        RECT 4.400 598.040 796.000 599.440 ;
        RECT 4.000 596.040 796.000 598.040 ;
        RECT 4.000 594.640 795.600 596.040 ;
        RECT 4.000 592.640 796.000 594.640 ;
        RECT 4.400 591.240 796.000 592.640 ;
        RECT 4.000 589.240 796.000 591.240 ;
        RECT 4.000 587.840 795.600 589.240 ;
        RECT 4.000 585.840 796.000 587.840 ;
        RECT 4.400 584.440 796.000 585.840 ;
        RECT 4.000 582.440 796.000 584.440 ;
        RECT 4.000 581.040 795.600 582.440 ;
        RECT 4.000 579.040 796.000 581.040 ;
        RECT 4.400 577.640 796.000 579.040 ;
        RECT 4.000 575.640 796.000 577.640 ;
        RECT 4.000 574.240 795.600 575.640 ;
        RECT 4.000 572.240 796.000 574.240 ;
        RECT 4.400 570.840 796.000 572.240 ;
        RECT 4.000 568.840 796.000 570.840 ;
        RECT 4.000 567.440 795.600 568.840 ;
        RECT 4.000 565.440 796.000 567.440 ;
        RECT 4.400 564.040 796.000 565.440 ;
        RECT 4.000 562.040 796.000 564.040 ;
        RECT 4.000 560.640 795.600 562.040 ;
        RECT 4.000 558.640 796.000 560.640 ;
        RECT 4.400 557.240 796.000 558.640 ;
        RECT 4.000 555.240 796.000 557.240 ;
        RECT 4.000 553.840 795.600 555.240 ;
        RECT 4.000 551.840 796.000 553.840 ;
        RECT 4.400 550.440 796.000 551.840 ;
        RECT 4.000 548.440 796.000 550.440 ;
        RECT 4.000 547.040 795.600 548.440 ;
        RECT 4.000 545.040 796.000 547.040 ;
        RECT 4.400 543.640 796.000 545.040 ;
        RECT 4.000 541.640 796.000 543.640 ;
        RECT 4.000 540.240 795.600 541.640 ;
        RECT 4.000 538.240 796.000 540.240 ;
        RECT 4.400 536.840 796.000 538.240 ;
        RECT 4.000 534.840 796.000 536.840 ;
        RECT 4.000 533.440 795.600 534.840 ;
        RECT 4.000 531.440 796.000 533.440 ;
        RECT 4.400 530.040 796.000 531.440 ;
        RECT 4.000 528.040 796.000 530.040 ;
        RECT 4.000 526.640 795.600 528.040 ;
        RECT 4.000 524.640 796.000 526.640 ;
        RECT 4.400 523.240 796.000 524.640 ;
        RECT 4.000 521.240 796.000 523.240 ;
        RECT 4.000 519.840 795.600 521.240 ;
        RECT 4.000 517.840 796.000 519.840 ;
        RECT 4.400 516.440 796.000 517.840 ;
        RECT 4.000 514.440 796.000 516.440 ;
        RECT 4.000 513.040 795.600 514.440 ;
        RECT 4.000 511.040 796.000 513.040 ;
        RECT 4.400 509.640 796.000 511.040 ;
        RECT 4.000 507.640 796.000 509.640 ;
        RECT 4.000 506.240 795.600 507.640 ;
        RECT 4.000 504.240 796.000 506.240 ;
        RECT 4.400 502.840 796.000 504.240 ;
        RECT 4.000 500.840 796.000 502.840 ;
        RECT 4.000 499.440 795.600 500.840 ;
        RECT 4.000 497.440 796.000 499.440 ;
        RECT 4.400 496.040 796.000 497.440 ;
        RECT 4.000 494.040 796.000 496.040 ;
        RECT 4.000 492.640 795.600 494.040 ;
        RECT 4.000 490.640 796.000 492.640 ;
        RECT 4.400 489.240 796.000 490.640 ;
        RECT 4.000 487.240 796.000 489.240 ;
        RECT 4.000 485.840 795.600 487.240 ;
        RECT 4.000 483.840 796.000 485.840 ;
        RECT 4.400 482.440 796.000 483.840 ;
        RECT 4.000 480.440 796.000 482.440 ;
        RECT 4.000 479.040 795.600 480.440 ;
        RECT 4.000 477.040 796.000 479.040 ;
        RECT 4.400 475.640 796.000 477.040 ;
        RECT 4.000 473.640 796.000 475.640 ;
        RECT 4.000 472.240 795.600 473.640 ;
        RECT 4.000 470.240 796.000 472.240 ;
        RECT 4.400 468.840 796.000 470.240 ;
        RECT 4.000 466.840 796.000 468.840 ;
        RECT 4.000 465.440 795.600 466.840 ;
        RECT 4.000 463.440 796.000 465.440 ;
        RECT 4.400 462.040 796.000 463.440 ;
        RECT 4.000 460.040 796.000 462.040 ;
        RECT 4.000 458.640 795.600 460.040 ;
        RECT 4.000 456.640 796.000 458.640 ;
        RECT 4.400 455.240 796.000 456.640 ;
        RECT 4.000 453.240 796.000 455.240 ;
        RECT 4.000 451.840 795.600 453.240 ;
        RECT 4.000 449.840 796.000 451.840 ;
        RECT 4.400 448.440 796.000 449.840 ;
        RECT 4.000 446.440 796.000 448.440 ;
        RECT 4.000 445.040 795.600 446.440 ;
        RECT 4.000 443.040 796.000 445.040 ;
        RECT 4.400 441.640 796.000 443.040 ;
        RECT 4.000 439.640 796.000 441.640 ;
        RECT 4.000 438.240 795.600 439.640 ;
        RECT 4.000 436.240 796.000 438.240 ;
        RECT 4.400 434.840 796.000 436.240 ;
        RECT 4.000 432.840 796.000 434.840 ;
        RECT 4.000 431.440 795.600 432.840 ;
        RECT 4.000 429.440 796.000 431.440 ;
        RECT 4.400 428.040 796.000 429.440 ;
        RECT 4.000 426.040 796.000 428.040 ;
        RECT 4.000 424.640 795.600 426.040 ;
        RECT 4.000 422.640 796.000 424.640 ;
        RECT 4.400 421.240 796.000 422.640 ;
        RECT 4.000 419.240 796.000 421.240 ;
        RECT 4.000 417.840 795.600 419.240 ;
        RECT 4.000 415.840 796.000 417.840 ;
        RECT 4.400 414.440 796.000 415.840 ;
        RECT 4.000 412.440 796.000 414.440 ;
        RECT 4.000 411.040 795.600 412.440 ;
        RECT 4.000 409.040 796.000 411.040 ;
        RECT 4.400 407.640 796.000 409.040 ;
        RECT 4.000 405.640 796.000 407.640 ;
        RECT 4.400 404.240 795.600 405.640 ;
        RECT 4.000 398.840 796.000 404.240 ;
        RECT 4.400 397.440 795.600 398.840 ;
        RECT 4.000 392.040 796.000 397.440 ;
        RECT 4.400 390.640 795.600 392.040 ;
        RECT 4.000 385.240 796.000 390.640 ;
        RECT 4.400 383.840 795.600 385.240 ;
        RECT 4.000 378.440 796.000 383.840 ;
        RECT 4.400 377.040 795.600 378.440 ;
        RECT 4.000 375.040 796.000 377.040 ;
        RECT 4.000 373.640 795.600 375.040 ;
        RECT 4.000 371.640 796.000 373.640 ;
        RECT 4.400 370.240 796.000 371.640 ;
        RECT 4.000 368.240 796.000 370.240 ;
        RECT 4.000 366.840 795.600 368.240 ;
        RECT 4.000 364.840 796.000 366.840 ;
        RECT 4.400 363.440 796.000 364.840 ;
        RECT 4.000 361.440 796.000 363.440 ;
        RECT 4.000 360.040 795.600 361.440 ;
        RECT 4.000 358.040 796.000 360.040 ;
        RECT 4.400 356.640 796.000 358.040 ;
        RECT 4.000 354.640 796.000 356.640 ;
        RECT 4.000 353.240 795.600 354.640 ;
        RECT 4.000 351.240 796.000 353.240 ;
        RECT 4.400 349.840 796.000 351.240 ;
        RECT 4.000 347.840 796.000 349.840 ;
        RECT 4.000 346.440 795.600 347.840 ;
        RECT 4.000 344.440 796.000 346.440 ;
        RECT 4.400 343.040 796.000 344.440 ;
        RECT 4.000 341.040 796.000 343.040 ;
        RECT 4.000 339.640 795.600 341.040 ;
        RECT 4.000 337.640 796.000 339.640 ;
        RECT 4.400 336.240 796.000 337.640 ;
        RECT 4.000 334.240 796.000 336.240 ;
        RECT 4.000 332.840 795.600 334.240 ;
        RECT 4.000 330.840 796.000 332.840 ;
        RECT 4.400 329.440 796.000 330.840 ;
        RECT 4.000 327.440 796.000 329.440 ;
        RECT 4.000 326.040 795.600 327.440 ;
        RECT 4.000 324.040 796.000 326.040 ;
        RECT 4.400 322.640 796.000 324.040 ;
        RECT 4.000 320.640 796.000 322.640 ;
        RECT 4.000 319.240 795.600 320.640 ;
        RECT 4.000 317.240 796.000 319.240 ;
        RECT 4.400 315.840 796.000 317.240 ;
        RECT 4.000 313.840 796.000 315.840 ;
        RECT 4.000 312.440 795.600 313.840 ;
        RECT 4.000 310.440 796.000 312.440 ;
        RECT 4.400 309.040 796.000 310.440 ;
        RECT 4.000 307.040 796.000 309.040 ;
        RECT 4.000 305.640 795.600 307.040 ;
        RECT 4.000 303.640 796.000 305.640 ;
        RECT 4.400 302.240 796.000 303.640 ;
        RECT 4.000 300.240 796.000 302.240 ;
        RECT 4.000 298.840 795.600 300.240 ;
        RECT 4.000 296.840 796.000 298.840 ;
        RECT 4.400 295.440 796.000 296.840 ;
        RECT 4.000 293.440 796.000 295.440 ;
        RECT 4.000 292.040 795.600 293.440 ;
        RECT 4.000 290.040 796.000 292.040 ;
        RECT 4.400 288.640 796.000 290.040 ;
        RECT 4.000 286.640 796.000 288.640 ;
        RECT 4.000 285.240 795.600 286.640 ;
        RECT 4.000 283.240 796.000 285.240 ;
        RECT 4.400 281.840 796.000 283.240 ;
        RECT 4.000 279.840 796.000 281.840 ;
        RECT 4.000 278.440 795.600 279.840 ;
        RECT 4.000 276.440 796.000 278.440 ;
        RECT 4.400 275.040 796.000 276.440 ;
        RECT 4.000 273.040 796.000 275.040 ;
        RECT 4.000 271.640 795.600 273.040 ;
        RECT 4.000 269.640 796.000 271.640 ;
        RECT 4.400 268.240 796.000 269.640 ;
        RECT 4.000 266.240 796.000 268.240 ;
        RECT 4.000 264.840 795.600 266.240 ;
        RECT 4.000 262.840 796.000 264.840 ;
        RECT 4.400 261.440 796.000 262.840 ;
        RECT 4.000 259.440 796.000 261.440 ;
        RECT 4.000 258.040 795.600 259.440 ;
        RECT 4.000 256.040 796.000 258.040 ;
        RECT 4.400 254.640 796.000 256.040 ;
        RECT 4.000 252.640 796.000 254.640 ;
        RECT 4.000 251.240 795.600 252.640 ;
        RECT 4.000 249.240 796.000 251.240 ;
        RECT 4.400 247.840 796.000 249.240 ;
        RECT 4.000 245.840 796.000 247.840 ;
        RECT 4.000 244.440 795.600 245.840 ;
        RECT 4.000 242.440 796.000 244.440 ;
        RECT 4.400 241.040 796.000 242.440 ;
        RECT 4.000 239.040 796.000 241.040 ;
        RECT 4.000 237.640 795.600 239.040 ;
        RECT 4.000 235.640 796.000 237.640 ;
        RECT 4.400 234.240 796.000 235.640 ;
        RECT 4.000 232.240 796.000 234.240 ;
        RECT 4.000 230.840 795.600 232.240 ;
        RECT 4.000 228.840 796.000 230.840 ;
        RECT 4.400 227.440 796.000 228.840 ;
        RECT 4.000 225.440 796.000 227.440 ;
        RECT 4.000 224.040 795.600 225.440 ;
        RECT 4.000 222.040 796.000 224.040 ;
        RECT 4.400 220.640 796.000 222.040 ;
        RECT 4.000 218.640 796.000 220.640 ;
        RECT 4.000 217.240 795.600 218.640 ;
        RECT 4.000 215.240 796.000 217.240 ;
        RECT 4.400 213.840 796.000 215.240 ;
        RECT 4.000 211.840 796.000 213.840 ;
        RECT 4.000 210.440 795.600 211.840 ;
        RECT 4.000 208.440 796.000 210.440 ;
        RECT 4.400 207.040 796.000 208.440 ;
        RECT 4.000 205.040 796.000 207.040 ;
        RECT 4.000 203.640 795.600 205.040 ;
        RECT 4.000 201.640 796.000 203.640 ;
        RECT 4.400 200.240 796.000 201.640 ;
        RECT 4.000 198.240 796.000 200.240 ;
        RECT 4.000 196.840 795.600 198.240 ;
        RECT 4.000 194.840 796.000 196.840 ;
        RECT 4.400 193.440 796.000 194.840 ;
        RECT 4.000 191.440 796.000 193.440 ;
        RECT 4.000 190.040 795.600 191.440 ;
        RECT 4.000 188.040 796.000 190.040 ;
        RECT 4.400 186.640 796.000 188.040 ;
        RECT 4.000 184.640 796.000 186.640 ;
        RECT 4.000 183.240 795.600 184.640 ;
        RECT 4.000 181.240 796.000 183.240 ;
        RECT 4.400 179.840 796.000 181.240 ;
        RECT 4.000 177.840 796.000 179.840 ;
        RECT 4.000 176.440 795.600 177.840 ;
        RECT 4.000 174.440 796.000 176.440 ;
        RECT 4.400 173.040 796.000 174.440 ;
        RECT 4.000 171.040 796.000 173.040 ;
        RECT 4.000 169.640 795.600 171.040 ;
        RECT 4.000 167.640 796.000 169.640 ;
        RECT 4.400 166.240 796.000 167.640 ;
        RECT 4.000 164.240 796.000 166.240 ;
        RECT 4.000 162.840 795.600 164.240 ;
        RECT 4.000 160.840 796.000 162.840 ;
        RECT 4.400 159.440 796.000 160.840 ;
        RECT 4.000 157.440 796.000 159.440 ;
        RECT 4.000 156.040 795.600 157.440 ;
        RECT 4.000 154.040 796.000 156.040 ;
        RECT 4.400 152.640 796.000 154.040 ;
        RECT 4.000 150.640 796.000 152.640 ;
        RECT 4.000 149.240 795.600 150.640 ;
        RECT 4.000 147.240 796.000 149.240 ;
        RECT 4.400 145.840 796.000 147.240 ;
        RECT 4.000 143.840 796.000 145.840 ;
        RECT 4.000 142.440 795.600 143.840 ;
        RECT 4.000 140.440 796.000 142.440 ;
        RECT 4.400 139.040 796.000 140.440 ;
        RECT 4.000 137.040 796.000 139.040 ;
        RECT 4.000 135.640 795.600 137.040 ;
        RECT 4.000 133.640 796.000 135.640 ;
        RECT 4.400 132.240 796.000 133.640 ;
        RECT 4.000 130.240 796.000 132.240 ;
        RECT 4.000 128.840 795.600 130.240 ;
        RECT 4.000 126.840 796.000 128.840 ;
        RECT 4.400 125.440 796.000 126.840 ;
        RECT 4.000 123.440 796.000 125.440 ;
        RECT 4.000 122.040 795.600 123.440 ;
        RECT 4.000 120.040 796.000 122.040 ;
        RECT 4.400 118.640 796.000 120.040 ;
        RECT 4.000 116.640 796.000 118.640 ;
        RECT 4.000 115.240 795.600 116.640 ;
        RECT 4.000 113.240 796.000 115.240 ;
        RECT 4.400 111.840 796.000 113.240 ;
        RECT 4.000 109.840 796.000 111.840 ;
        RECT 4.000 108.440 795.600 109.840 ;
        RECT 4.000 106.440 796.000 108.440 ;
        RECT 4.400 105.040 796.000 106.440 ;
        RECT 4.000 103.040 796.000 105.040 ;
        RECT 4.000 101.640 795.600 103.040 ;
        RECT 4.000 99.640 796.000 101.640 ;
        RECT 4.400 98.240 796.000 99.640 ;
        RECT 4.000 96.240 796.000 98.240 ;
        RECT 4.000 94.840 795.600 96.240 ;
        RECT 4.000 92.840 796.000 94.840 ;
        RECT 4.400 91.440 796.000 92.840 ;
        RECT 4.000 89.440 796.000 91.440 ;
        RECT 4.000 88.040 795.600 89.440 ;
        RECT 4.000 86.040 796.000 88.040 ;
        RECT 4.400 84.640 796.000 86.040 ;
        RECT 4.000 82.640 796.000 84.640 ;
        RECT 4.000 81.240 795.600 82.640 ;
        RECT 4.000 79.240 796.000 81.240 ;
        RECT 4.400 77.840 796.000 79.240 ;
        RECT 4.000 75.840 796.000 77.840 ;
        RECT 4.000 74.440 795.600 75.840 ;
        RECT 4.000 72.440 796.000 74.440 ;
        RECT 4.400 71.040 796.000 72.440 ;
        RECT 4.000 69.040 796.000 71.040 ;
        RECT 4.000 67.640 795.600 69.040 ;
        RECT 4.000 65.640 796.000 67.640 ;
        RECT 4.400 64.240 796.000 65.640 ;
        RECT 4.000 62.240 796.000 64.240 ;
        RECT 4.000 60.840 795.600 62.240 ;
        RECT 4.000 58.840 796.000 60.840 ;
        RECT 4.400 57.440 796.000 58.840 ;
        RECT 4.000 55.440 796.000 57.440 ;
        RECT 4.000 54.040 795.600 55.440 ;
        RECT 4.000 52.040 796.000 54.040 ;
        RECT 4.400 50.640 796.000 52.040 ;
        RECT 4.000 48.640 796.000 50.640 ;
        RECT 4.000 47.240 795.600 48.640 ;
        RECT 4.000 45.240 796.000 47.240 ;
        RECT 4.400 43.840 796.000 45.240 ;
        RECT 4.000 41.840 796.000 43.840 ;
        RECT 4.000 40.440 795.600 41.840 ;
        RECT 4.000 38.440 796.000 40.440 ;
        RECT 4.400 37.040 796.000 38.440 ;
        RECT 4.000 35.040 796.000 37.040 ;
        RECT 4.000 33.640 795.600 35.040 ;
        RECT 4.000 31.640 796.000 33.640 ;
        RECT 4.400 30.240 796.000 31.640 ;
        RECT 4.000 28.240 796.000 30.240 ;
        RECT 4.000 26.840 795.600 28.240 ;
        RECT 4.000 24.840 796.000 26.840 ;
        RECT 4.400 23.440 796.000 24.840 ;
        RECT 4.000 21.440 796.000 23.440 ;
        RECT 4.000 20.040 795.600 21.440 ;
        RECT 4.000 18.040 796.000 20.040 ;
        RECT 4.400 16.640 796.000 18.040 ;
        RECT 4.000 14.640 796.000 16.640 ;
        RECT 4.000 13.240 795.600 14.640 ;
        RECT 4.000 11.240 796.000 13.240 ;
        RECT 4.400 9.840 796.000 11.240 ;
        RECT 4.000 7.840 796.000 9.840 ;
        RECT 4.000 6.440 795.600 7.840 ;
        RECT 4.000 4.440 796.000 6.440 ;
        RECT 4.400 3.040 796.000 4.440 ;
        RECT 4.000 1.040 796.000 3.040 ;
        RECT 4.000 0.175 795.600 1.040 ;
      LAYER met4 ;
        RECT 319.535 413.615 327.840 1244.905 ;
        RECT 330.240 413.615 404.640 1244.905 ;
        RECT 407.040 413.615 428.425 1244.905 ;
  END
END user_proj_example
END LIBRARY

