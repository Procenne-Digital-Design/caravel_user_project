VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO trng_wb_wrapper
  CLASS BLOCK ;
  FOREIGN trng_wb_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 1000.000 ;
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 455.640 750.000 456.240 ;
    END
  END rst_i
  PIN trng_buffer_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 996.000 203.230 1000.000 ;
    END
  END trng_buffer_o[0]
  PIN trng_buffer_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END trng_buffer_o[10]
  PIN trng_buffer_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 996.000 415.750 1000.000 ;
    END
  END trng_buffer_o[11]
  PIN trng_buffer_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END trng_buffer_o[12]
  PIN trng_buffer_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END trng_buffer_o[13]
  PIN trng_buffer_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END trng_buffer_o[14]
  PIN trng_buffer_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END trng_buffer_o[15]
  PIN trng_buffer_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 996.000 174.250 1000.000 ;
    END
  END trng_buffer_o[16]
  PIN trng_buffer_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END trng_buffer_o[17]
  PIN trng_buffer_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END trng_buffer_o[18]
  PIN trng_buffer_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 996.000 657.250 1000.000 ;
    END
  END trng_buffer_o[19]
  PIN trng_buffer_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 71.440 750.000 72.040 ;
    END
  END trng_buffer_o[1]
  PIN trng_buffer_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 901.040 750.000 901.640 ;
    END
  END trng_buffer_o[20]
  PIN trng_buffer_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END trng_buffer_o[21]
  PIN trng_buffer_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 166.640 750.000 167.240 ;
    END
  END trng_buffer_o[22]
  PIN trng_buffer_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 836.440 750.000 837.040 ;
    END
  END trng_buffer_o[23]
  PIN trng_buffer_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 996.000 325.590 1000.000 ;
    END
  END trng_buffer_o[24]
  PIN trng_buffer_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 996.000 22.910 1000.000 ;
    END
  END trng_buffer_o[25]
  PIN trng_buffer_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 935.040 750.000 935.640 ;
    END
  END trng_buffer_o[26]
  PIN trng_buffer_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 996.000 113.070 1000.000 ;
    END
  END trng_buffer_o[27]
  PIN trng_buffer_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END trng_buffer_o[28]
  PIN trng_buffer_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 37.440 750.000 38.040 ;
    END
  END trng_buffer_o[29]
  PIN trng_buffer_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END trng_buffer_o[2]
  PIN trng_buffer_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 996.000 354.570 1000.000 ;
    END
  END trng_buffer_o[30]
  PIN trng_buffer_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END trng_buffer_o[31]
  PIN trng_buffer_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END trng_buffer_o[3]
  PIN trng_buffer_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 996.000 264.410 1000.000 ;
    END
  END trng_buffer_o[4]
  PIN trng_buffer_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 326.440 750.000 327.040 ;
    END
  END trng_buffer_o[5]
  PIN trng_buffer_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END trng_buffer_o[6]
  PIN trng_buffer_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END trng_buffer_o[7]
  PIN trng_buffer_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END trng_buffer_o[8]
  PIN trng_buffer_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 996.000 596.070 1000.000 ;
    END
  END trng_buffer_o[9]
  PIN trng_valid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END trng_valid_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 357.040 750.000 357.640 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 870.440 750.000 871.040 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 775.240 750.000 775.840 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 710.640 750.000 711.240 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 676.640 750.000 677.240 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 965.640 750.000 966.240 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 996.000 293.390 1000.000 ;
    END
  END wb_adr_i[8]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 550.840 750.000 551.440 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 581.440 750.000 582.040 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 996.000 142.050 1000.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 996.000 386.770 1000.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 996.000 689.450 1000.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 292.440 750.000 293.040 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 197.240 750.000 197.840 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 6.840 750.000 7.440 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 261.840 750.000 262.440 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 996.000 747.410 1000.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 391.040 750.000 391.640 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 996.000 80.870 1000.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 132.640 750.000 133.240 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 996.000 476.930 1000.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 102.040 750.000 102.640 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 615.440 750.000 616.040 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 421.640 750.000 422.240 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 486.240 750.000 486.840 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 741.240 750.000 741.840 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 805.840 750.000 806.440 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 996.000 235.430 1000.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 996.000 505.910 1000.000 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 996.000 628.270 1000.000 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 996.000 444.730 1000.000 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 996.000 718.430 1000.000 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 231.240 750.000 231.840 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 646.040 750.000 646.640 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 996.000 567.090 1000.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 996.000 538.110 1000.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 996.000 51.890 1000.000 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wb_dat_o[9]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 516.840 750.000 517.440 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 744.280 987.445 ;
      LAYER met1 ;
        RECT 0.070 10.640 749.730 987.600 ;
      LAYER met2 ;
        RECT 0.100 995.720 22.350 996.610 ;
        RECT 23.190 995.720 51.330 996.610 ;
        RECT 52.170 995.720 80.310 996.610 ;
        RECT 81.150 995.720 112.510 996.610 ;
        RECT 113.350 995.720 141.490 996.610 ;
        RECT 142.330 995.720 173.690 996.610 ;
        RECT 174.530 995.720 202.670 996.610 ;
        RECT 203.510 995.720 234.870 996.610 ;
        RECT 235.710 995.720 263.850 996.610 ;
        RECT 264.690 995.720 292.830 996.610 ;
        RECT 293.670 995.720 325.030 996.610 ;
        RECT 325.870 995.720 354.010 996.610 ;
        RECT 354.850 995.720 386.210 996.610 ;
        RECT 387.050 995.720 415.190 996.610 ;
        RECT 416.030 995.720 444.170 996.610 ;
        RECT 445.010 995.720 476.370 996.610 ;
        RECT 477.210 995.720 505.350 996.610 ;
        RECT 506.190 995.720 537.550 996.610 ;
        RECT 538.390 995.720 566.530 996.610 ;
        RECT 567.370 995.720 595.510 996.610 ;
        RECT 596.350 995.720 627.710 996.610 ;
        RECT 628.550 995.720 656.690 996.610 ;
        RECT 657.530 995.720 688.890 996.610 ;
        RECT 689.730 995.720 717.870 996.610 ;
        RECT 718.710 995.720 746.850 996.610 ;
        RECT 747.690 995.720 749.700 996.610 ;
        RECT 0.100 4.280 749.700 995.720 ;
        RECT 0.650 4.000 28.790 4.280 ;
        RECT 29.630 4.000 57.770 4.280 ;
        RECT 58.610 4.000 89.970 4.280 ;
        RECT 90.810 4.000 118.950 4.280 ;
        RECT 119.790 4.000 151.150 4.280 ;
        RECT 151.990 4.000 180.130 4.280 ;
        RECT 180.970 4.000 209.110 4.280 ;
        RECT 209.950 4.000 241.310 4.280 ;
        RECT 242.150 4.000 270.290 4.280 ;
        RECT 271.130 4.000 302.490 4.280 ;
        RECT 303.330 4.000 331.470 4.280 ;
        RECT 332.310 4.000 360.450 4.280 ;
        RECT 361.290 4.000 392.650 4.280 ;
        RECT 393.490 4.000 421.630 4.280 ;
        RECT 422.470 4.000 453.830 4.280 ;
        RECT 454.670 4.000 482.810 4.280 ;
        RECT 483.650 4.000 511.790 4.280 ;
        RECT 512.630 4.000 543.990 4.280 ;
        RECT 544.830 4.000 572.970 4.280 ;
        RECT 573.810 4.000 605.170 4.280 ;
        RECT 606.010 4.000 634.150 4.280 ;
        RECT 634.990 4.000 666.350 4.280 ;
        RECT 667.190 4.000 695.330 4.280 ;
        RECT 696.170 4.000 724.310 4.280 ;
        RECT 725.150 4.000 749.700 4.280 ;
      LAYER met3 ;
        RECT 4.400 989.040 748.815 989.905 ;
        RECT 4.000 966.640 748.815 989.040 ;
        RECT 4.000 965.240 745.600 966.640 ;
        RECT 4.000 959.840 748.815 965.240 ;
        RECT 4.400 958.440 748.815 959.840 ;
        RECT 4.000 936.040 748.815 958.440 ;
        RECT 4.000 934.640 745.600 936.040 ;
        RECT 4.000 925.840 748.815 934.640 ;
        RECT 4.400 924.440 748.815 925.840 ;
        RECT 4.000 902.040 748.815 924.440 ;
        RECT 4.000 900.640 745.600 902.040 ;
        RECT 4.000 895.240 748.815 900.640 ;
        RECT 4.400 893.840 748.815 895.240 ;
        RECT 4.000 871.440 748.815 893.840 ;
        RECT 4.000 870.040 745.600 871.440 ;
        RECT 4.000 864.640 748.815 870.040 ;
        RECT 4.400 863.240 748.815 864.640 ;
        RECT 4.000 837.440 748.815 863.240 ;
        RECT 4.000 836.040 745.600 837.440 ;
        RECT 4.000 830.640 748.815 836.040 ;
        RECT 4.400 829.240 748.815 830.640 ;
        RECT 4.000 806.840 748.815 829.240 ;
        RECT 4.000 805.440 745.600 806.840 ;
        RECT 4.000 800.040 748.815 805.440 ;
        RECT 4.400 798.640 748.815 800.040 ;
        RECT 4.000 776.240 748.815 798.640 ;
        RECT 4.000 774.840 745.600 776.240 ;
        RECT 4.000 766.040 748.815 774.840 ;
        RECT 4.400 764.640 748.815 766.040 ;
        RECT 4.000 742.240 748.815 764.640 ;
        RECT 4.000 740.840 745.600 742.240 ;
        RECT 4.000 735.440 748.815 740.840 ;
        RECT 4.400 734.040 748.815 735.440 ;
        RECT 4.000 711.640 748.815 734.040 ;
        RECT 4.000 710.240 745.600 711.640 ;
        RECT 4.000 704.840 748.815 710.240 ;
        RECT 4.400 703.440 748.815 704.840 ;
        RECT 4.000 677.640 748.815 703.440 ;
        RECT 4.000 676.240 745.600 677.640 ;
        RECT 4.000 670.840 748.815 676.240 ;
        RECT 4.400 669.440 748.815 670.840 ;
        RECT 4.000 647.040 748.815 669.440 ;
        RECT 4.000 645.640 745.600 647.040 ;
        RECT 4.000 640.240 748.815 645.640 ;
        RECT 4.400 638.840 748.815 640.240 ;
        RECT 4.000 616.440 748.815 638.840 ;
        RECT 4.000 615.040 745.600 616.440 ;
        RECT 4.000 606.240 748.815 615.040 ;
        RECT 4.400 604.840 748.815 606.240 ;
        RECT 4.000 582.440 748.815 604.840 ;
        RECT 4.000 581.040 745.600 582.440 ;
        RECT 4.000 575.640 748.815 581.040 ;
        RECT 4.400 574.240 748.815 575.640 ;
        RECT 4.000 551.840 748.815 574.240 ;
        RECT 4.000 550.440 745.600 551.840 ;
        RECT 4.000 541.640 748.815 550.440 ;
        RECT 4.400 540.240 748.815 541.640 ;
        RECT 4.000 517.840 748.815 540.240 ;
        RECT 4.000 516.440 745.600 517.840 ;
        RECT 4.000 511.040 748.815 516.440 ;
        RECT 4.400 509.640 748.815 511.040 ;
        RECT 4.000 487.240 748.815 509.640 ;
        RECT 4.000 485.840 745.600 487.240 ;
        RECT 4.000 480.440 748.815 485.840 ;
        RECT 4.400 479.040 748.815 480.440 ;
        RECT 4.000 456.640 748.815 479.040 ;
        RECT 4.000 455.240 745.600 456.640 ;
        RECT 4.000 446.440 748.815 455.240 ;
        RECT 4.400 445.040 748.815 446.440 ;
        RECT 4.000 422.640 748.815 445.040 ;
        RECT 4.000 421.240 745.600 422.640 ;
        RECT 4.000 415.840 748.815 421.240 ;
        RECT 4.400 414.440 748.815 415.840 ;
        RECT 4.000 392.040 748.815 414.440 ;
        RECT 4.000 390.640 745.600 392.040 ;
        RECT 4.000 381.840 748.815 390.640 ;
        RECT 4.400 380.440 748.815 381.840 ;
        RECT 4.000 358.040 748.815 380.440 ;
        RECT 4.000 356.640 745.600 358.040 ;
        RECT 4.000 351.240 748.815 356.640 ;
        RECT 4.400 349.840 748.815 351.240 ;
        RECT 4.000 327.440 748.815 349.840 ;
        RECT 4.000 326.040 745.600 327.440 ;
        RECT 4.000 320.640 748.815 326.040 ;
        RECT 4.400 319.240 748.815 320.640 ;
        RECT 4.000 293.440 748.815 319.240 ;
        RECT 4.000 292.040 745.600 293.440 ;
        RECT 4.000 286.640 748.815 292.040 ;
        RECT 4.400 285.240 748.815 286.640 ;
        RECT 4.000 262.840 748.815 285.240 ;
        RECT 4.000 261.440 745.600 262.840 ;
        RECT 4.000 256.040 748.815 261.440 ;
        RECT 4.400 254.640 748.815 256.040 ;
        RECT 4.000 232.240 748.815 254.640 ;
        RECT 4.000 230.840 745.600 232.240 ;
        RECT 4.000 222.040 748.815 230.840 ;
        RECT 4.400 220.640 748.815 222.040 ;
        RECT 4.000 198.240 748.815 220.640 ;
        RECT 4.000 196.840 745.600 198.240 ;
        RECT 4.000 191.440 748.815 196.840 ;
        RECT 4.400 190.040 748.815 191.440 ;
        RECT 4.000 167.640 748.815 190.040 ;
        RECT 4.000 166.240 745.600 167.640 ;
        RECT 4.000 160.840 748.815 166.240 ;
        RECT 4.400 159.440 748.815 160.840 ;
        RECT 4.000 133.640 748.815 159.440 ;
        RECT 4.000 132.240 745.600 133.640 ;
        RECT 4.000 126.840 748.815 132.240 ;
        RECT 4.400 125.440 748.815 126.840 ;
        RECT 4.000 103.040 748.815 125.440 ;
        RECT 4.000 101.640 745.600 103.040 ;
        RECT 4.000 96.240 748.815 101.640 ;
        RECT 4.400 94.840 748.815 96.240 ;
        RECT 4.000 72.440 748.815 94.840 ;
        RECT 4.000 71.040 745.600 72.440 ;
        RECT 4.000 62.240 748.815 71.040 ;
        RECT 4.400 60.840 748.815 62.240 ;
        RECT 4.000 38.440 748.815 60.840 ;
        RECT 4.000 37.040 745.600 38.440 ;
        RECT 4.000 31.640 748.815 37.040 ;
        RECT 4.400 30.240 748.815 31.640 ;
        RECT 4.000 10.715 748.815 30.240 ;
      LAYER met4 ;
        RECT 495.255 351.735 558.240 760.065 ;
        RECT 560.640 351.735 635.040 760.065 ;
        RECT 637.440 351.735 711.840 760.065 ;
        RECT 714.240 351.735 748.585 760.065 ;
  END
END trng_wb_wrapper
END LIBRARY

