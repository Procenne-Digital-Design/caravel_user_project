VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_interconnect
  CLASS BLOCK ;
  FOREIGN wb_interconnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 1200.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1196.000 193.570 1200.000 ;
    END
  END clk_i
  PIN m0_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1173.040 400.000 1173.640 ;
    END
  END m0_wb_ack_o
  PIN m0_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END m0_wb_adr_i[0]
  PIN m0_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 860.240 400.000 860.840 ;
    END
  END m0_wb_adr_i[10]
  PIN m0_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END m0_wb_adr_i[11]
  PIN m0_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.040 400.000 204.640 ;
    END
  END m0_wb_adr_i[12]
  PIN m0_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END m0_wb_adr_i[13]
  PIN m0_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END m0_wb_adr_i[14]
  PIN m0_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 544.040 400.000 544.640 ;
    END
  END m0_wb_adr_i[15]
  PIN m0_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1196.000 251.530 1200.000 ;
    END
  END m0_wb_adr_i[16]
  PIN m0_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END m0_wb_adr_i[17]
  PIN m0_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END m0_wb_adr_i[18]
  PIN m0_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1115.240 400.000 1115.840 ;
    END
  END m0_wb_adr_i[19]
  PIN m0_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END m0_wb_adr_i[1]
  PIN m0_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 737.840 400.000 738.440 ;
    END
  END m0_wb_adr_i[20]
  PIN m0_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 676.640 400.000 677.240 ;
    END
  END m0_wb_adr_i[21]
  PIN m0_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1064.240 400.000 1064.840 ;
    END
  END m0_wb_adr_i[22]
  PIN m0_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END m0_wb_adr_i[23]
  PIN m0_wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END m0_wb_adr_i[24]
  PIN m0_wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 506.640 400.000 507.240 ;
    END
  END m0_wb_adr_i[25]
  PIN m0_wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1196.000 10.030 1200.000 ;
    END
  END m0_wb_adr_i[26]
  PIN m0_wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 387.640 400.000 388.240 ;
    END
  END m0_wb_adr_i[27]
  PIN m0_wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1196.000 309.490 1200.000 ;
    END
  END m0_wb_adr_i[28]
  PIN m0_wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END m0_wb_adr_i[29]
  PIN m0_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 275.440 400.000 276.040 ;
    END
  END m0_wb_adr_i[2]
  PIN m0_wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END m0_wb_adr_i[30]
  PIN m0_wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 166.640 400.000 167.240 ;
    END
  END m0_wb_adr_i[31]
  PIN m0_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 241.440 400.000 242.040 ;
    END
  END m0_wb_adr_i[3]
  PIN m0_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 809.240 400.000 809.840 ;
    END
  END m0_wb_adr_i[4]
  PIN m0_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1077.840 400.000 1078.440 ;
    END
  END m0_wb_adr_i[5]
  PIN m0_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END m0_wb_adr_i[6]
  PIN m0_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 326.440 400.000 327.040 ;
    END
  END m0_wb_adr_i[7]
  PIN m0_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END m0_wb_adr_i[8]
  PIN m0_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 799.040 400.000 799.640 ;
    END
  END m0_wb_adr_i[9]
  PIN m0_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.040 400.000 119.640 ;
    END
  END m0_wb_cyc_i
  PIN m0_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END m0_wb_dat_i[0]
  PIN m0_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END m0_wb_dat_i[10]
  PIN m0_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 71.440 400.000 72.040 ;
    END
  END m0_wb_dat_i[11]
  PIN m0_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END m0_wb_dat_i[12]
  PIN m0_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 979.240 400.000 979.840 ;
    END
  END m0_wb_dat_i[13]
  PIN m0_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END m0_wb_dat_i[14]
  PIN m0_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END m0_wb_dat_i[15]
  PIN m0_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END m0_wb_dat_i[16]
  PIN m0_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1196.000 367.450 1200.000 ;
    END
  END m0_wb_dat_i[17]
  PIN m0_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END m0_wb_dat_i[18]
  PIN m0_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END m0_wb_dat_i[19]
  PIN m0_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END m0_wb_dat_i[1]
  PIN m0_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.840 400.000 398.440 ;
    END
  END m0_wb_dat_i[20]
  PIN m0_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END m0_wb_dat_i[21]
  PIN m0_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 496.440 400.000 497.040 ;
    END
  END m0_wb_dat_i[22]
  PIN m0_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END m0_wb_dat_i[23]
  PIN m0_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END m0_wb_dat_i[24]
  PIN m0_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 629.040 400.000 629.640 ;
    END
  END m0_wb_dat_i[25]
  PIN m0_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 918.040 400.000 918.640 ;
    END
  END m0_wb_dat_i[26]
  PIN m0_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END m0_wb_dat_i[27]
  PIN m0_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END m0_wb_dat_i[28]
  PIN m0_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1196.000 67.990 1200.000 ;
    END
  END m0_wb_dat_i[29]
  PIN m0_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END m0_wb_dat_i[2]
  PIN m0_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END m0_wb_dat_i[30]
  PIN m0_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END m0_wb_dat_i[31]
  PIN m0_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END m0_wb_dat_i[3]
  PIN m0_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1196.000 113.070 1200.000 ;
    END
  END m0_wb_dat_i[4]
  PIN m0_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END m0_wb_dat_i[5]
  PIN m0_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1196.000 90.530 1200.000 ;
    END
  END m0_wb_dat_i[6]
  PIN m0_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1196.000 183.910 1200.000 ;
    END
  END m0_wb_dat_i[7]
  PIN m0_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 1196.000 125.950 1200.000 ;
    END
  END m0_wb_dat_i[8]
  PIN m0_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 302.640 400.000 303.240 ;
    END
  END m0_wb_dat_i[9]
  PIN m0_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1149.240 400.000 1149.840 ;
    END
  END m0_wb_dat_o[0]
  PIN m0_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END m0_wb_dat_o[10]
  PIN m0_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END m0_wb_dat_o[11]
  PIN m0_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 459.040 400.000 459.640 ;
    END
  END m0_wb_dat_o[12]
  PIN m0_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END m0_wb_dat_o[13]
  PIN m0_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 945.240 400.000 945.840 ;
    END
  END m0_wb_dat_o[14]
  PIN m0_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1186.640 4.000 1187.240 ;
    END
  END m0_wb_dat_o[15]
  PIN m0_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 217.640 400.000 218.240 ;
    END
  END m0_wb_dat_o[16]
  PIN m0_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END m0_wb_dat_o[17]
  PIN m0_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END m0_wb_dat_o[18]
  PIN m0_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.040 400.000 34.640 ;
    END
  END m0_wb_dat_o[19]
  PIN m0_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END m0_wb_dat_o[1]
  PIN m0_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 605.240 400.000 605.840 ;
    END
  END m0_wb_dat_o[20]
  PIN m0_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 1196.000 389.990 1200.000 ;
    END
  END m0_wb_dat_o[21]
  PIN m0_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END m0_wb_dat_o[22]
  PIN m0_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END m0_wb_dat_o[23]
  PIN m0_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 336.640 400.000 337.240 ;
    END
  END m0_wb_dat_o[24]
  PIN m0_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END m0_wb_dat_o[25]
  PIN m0_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.840 400.000 313.440 ;
    END
  END m0_wb_dat_o[26]
  PIN m0_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1003.040 400.000 1003.640 ;
    END
  END m0_wb_dat_o[27]
  PIN m0_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END m0_wb_dat_o[28]
  PIN m0_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 822.840 400.000 823.440 ;
    END
  END m0_wb_dat_o[29]
  PIN m0_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 81.640 400.000 82.240 ;
    END
  END m0_wb_dat_o[2]
  PIN m0_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END m0_wb_dat_o[30]
  PIN m0_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END m0_wb_dat_o[31]
  PIN m0_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 1196.000 241.870 1200.000 ;
    END
  END m0_wb_dat_o[3]
  PIN m0_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END m0_wb_dat_o[4]
  PIN m0_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 251.640 400.000 252.240 ;
    END
  END m0_wb_dat_o[5]
  PIN m0_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END m0_wb_dat_o[6]
  PIN m0_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1196.000 22.910 1200.000 ;
    END
  END m0_wb_dat_o[7]
  PIN m0_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 884.040 400.000 884.640 ;
    END
  END m0_wb_dat_o[8]
  PIN m0_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 846.640 400.000 847.240 ;
    END
  END m0_wb_dat_o[9]
  PIN m0_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1196.000 0.370 1200.000 ;
    END
  END m0_wb_sel_i[0]
  PIN m0_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1196.000 32.570 1200.000 ;
    END
  END m0_wb_sel_i[1]
  PIN m0_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END m0_wb_sel_i[2]
  PIN m0_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END m0_wb_sel_i[3]
  PIN m0_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END m0_wb_stb_i
  PIN m0_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.840 400.000 143.440 ;
    END
  END m0_wb_we_i
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END rst_n
  PIN s0_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END s0_wb_ack_i
  PIN s0_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 700.440 400.000 701.040 ;
    END
  END s0_wb_adr_o[0]
  PIN s0_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1040.440 400.000 1041.040 ;
    END
  END s0_wb_adr_o[1]
  PIN s0_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END s0_wb_adr_o[2]
  PIN s0_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 445.440 400.000 446.040 ;
    END
  END s0_wb_adr_o[3]
  PIN s0_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END s0_wb_adr_o[4]
  PIN s0_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 833.040 400.000 833.640 ;
    END
  END s0_wb_adr_o[5]
  PIN s0_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END s0_wb_adr_o[6]
  PIN s0_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 411.440 400.000 412.040 ;
    END
  END s0_wb_adr_o[7]
  PIN s0_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 652.840 400.000 653.440 ;
    END
  END s0_wb_adr_o[8]
  PIN s0_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END s0_wb_cyc_o
  PIN s0_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 615.440 400.000 616.040 ;
    END
  END s0_wb_dat_i[0]
  PIN s0_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END s0_wb_dat_i[10]
  PIN s0_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 1196.000 354.570 1200.000 ;
    END
  END s0_wb_dat_i[11]
  PIN s0_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END s0_wb_dat_i[12]
  PIN s0_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 775.240 400.000 775.840 ;
    END
  END s0_wb_dat_i[13]
  PIN s0_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END s0_wb_dat_i[14]
  PIN s0_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END s0_wb_dat_i[15]
  PIN s0_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 10.240 400.000 10.840 ;
    END
  END s0_wb_dat_i[16]
  PIN s0_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END s0_wb_dat_i[17]
  PIN s0_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 1196.000 322.370 1200.000 ;
    END
  END s0_wb_dat_i[18]
  PIN s0_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END s0_wb_dat_i[19]
  PIN s0_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END s0_wb_dat_i[1]
  PIN s0_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END s0_wb_dat_i[20]
  PIN s0_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END s0_wb_dat_i[21]
  PIN s0_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END s0_wb_dat_i[22]
  PIN s0_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END s0_wb_dat_i[23]
  PIN s0_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 870.440 400.000 871.040 ;
    END
  END s0_wb_dat_i[24]
  PIN s0_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END s0_wb_dat_i[25]
  PIN s0_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END s0_wb_dat_i[26]
  PIN s0_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 20.440 400.000 21.040 ;
    END
  END s0_wb_dat_i[27]
  PIN s0_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1196.000 55.110 1200.000 ;
    END
  END s0_wb_dat_i[28]
  PIN s0_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END s0_wb_dat_i[29]
  PIN s0_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 1196.000 216.110 1200.000 ;
    END
  END s0_wb_dat_i[2]
  PIN s0_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 1196.000 377.110 1200.000 ;
    END
  END s0_wb_dat_i[30]
  PIN s0_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END s0_wb_dat_i[31]
  PIN s0_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END s0_wb_dat_i[3]
  PIN s0_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1016.640 400.000 1017.240 ;
    END
  END s0_wb_dat_i[4]
  PIN s0_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 520.240 400.000 520.840 ;
    END
  END s0_wb_dat_i[5]
  PIN s0_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 47.640 400.000 48.240 ;
    END
  END s0_wb_dat_i[6]
  PIN s0_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 894.240 400.000 894.840 ;
    END
  END s0_wb_dat_i[7]
  PIN s0_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.240 400.000 265.840 ;
    END
  END s0_wb_dat_i[8]
  PIN s0_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END s0_wb_dat_i[9]
  PIN s0_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END s0_wb_dat_o[0]
  PIN s0_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1196.000 135.610 1200.000 ;
    END
  END s0_wb_dat_o[10]
  PIN s0_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END s0_wb_dat_o[11]
  PIN s0_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 530.440 400.000 531.040 ;
    END
  END s0_wb_dat_o[12]
  PIN s0_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END s0_wb_dat_o[13]
  PIN s0_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 639.240 400.000 639.840 ;
    END
  END s0_wb_dat_o[14]
  PIN s0_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END s0_wb_dat_o[15]
  PIN s0_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END s0_wb_dat_o[16]
  PIN s0_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 1196.000 274.070 1200.000 ;
    END
  END s0_wb_dat_o[17]
  PIN s0_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END s0_wb_dat_o[18]
  PIN s0_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 724.240 400.000 724.840 ;
    END
  END s0_wb_dat_o[19]
  PIN s0_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 1196.000 228.990 1200.000 ;
    END
  END s0_wb_dat_o[1]
  PIN s0_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1196.000 286.950 1200.000 ;
    END
  END s0_wb_dat_o[20]
  PIN s0_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 350.240 400.000 350.840 ;
    END
  END s0_wb_dat_o[21]
  PIN s0_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END s0_wb_dat_o[22]
  PIN s0_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END s0_wb_dat_o[23]
  PIN s0_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1125.440 400.000 1126.040 ;
    END
  END s0_wb_dat_o[24]
  PIN s0_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END s0_wb_dat_o[25]
  PIN s0_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END s0_wb_dat_o[26]
  PIN s0_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END s0_wb_dat_o[27]
  PIN s0_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END s0_wb_dat_o[28]
  PIN s0_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 751.440 400.000 752.040 ;
    END
  END s0_wb_dat_o[29]
  PIN s0_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 714.040 400.000 714.640 ;
    END
  END s0_wb_dat_o[2]
  PIN s0_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END s0_wb_dat_o[30]
  PIN s0_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END s0_wb_dat_o[31]
  PIN s0_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 469.240 400.000 469.840 ;
    END
  END s0_wb_dat_o[3]
  PIN s0_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.840 400.000 228.440 ;
    END
  END s0_wb_dat_o[4]
  PIN s0_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1186.640 400.000 1187.240 ;
    END
  END s0_wb_dat_o[5]
  PIN s0_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END s0_wb_dat_o[6]
  PIN s0_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END s0_wb_dat_o[7]
  PIN s0_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END s0_wb_dat_o[8]
  PIN s0_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 421.640 400.000 422.240 ;
    END
  END s0_wb_dat_o[9]
  PIN s0_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1196.000 45.450 1200.000 ;
    END
  END s0_wb_sel_o[0]
  PIN s0_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END s0_wb_sel_o[1]
  PIN s0_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END s0_wb_sel_o[2]
  PIN s0_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1196.000 171.030 1200.000 ;
    END
  END s0_wb_sel_o[3]
  PIN s0_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END s0_wb_stb_o
  PIN s0_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 955.440 400.000 956.040 ;
    END
  END s0_wb_we_o
  PIN s1_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END s1_wb_ack_i
  PIN s1_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1139.040 400.000 1139.640 ;
    END
  END s1_wb_adr_o[0]
  PIN s1_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 581.440 400.000 582.040 ;
    END
  END s1_wb_adr_o[1]
  PIN s1_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 132.640 400.000 133.240 ;
    END
  END s1_wb_adr_o[2]
  PIN s1_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1162.840 400.000 1163.440 ;
    END
  END s1_wb_adr_o[3]
  PIN s1_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 105.440 400.000 106.040 ;
    END
  END s1_wb_adr_o[4]
  PIN s1_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END s1_wb_adr_o[5]
  PIN s1_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END s1_wb_adr_o[6]
  PIN s1_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.040 400.000 289.640 ;
    END
  END s1_wb_adr_o[7]
  PIN s1_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 482.840 400.000 483.440 ;
    END
  END s1_wb_adr_o[8]
  PIN s1_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1196.000 103.410 1200.000 ;
    END
  END s1_wb_cyc_o
  PIN s1_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 931.640 400.000 932.240 ;
    END
  END s1_wb_dat_i[0]
  PIN s1_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END s1_wb_dat_i[10]
  PIN s1_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END s1_wb_dat_i[11]
  PIN s1_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END s1_wb_dat_i[12]
  PIN s1_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END s1_wb_dat_i[13]
  PIN s1_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END s1_wb_dat_i[14]
  PIN s1_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 690.240 400.000 690.840 ;
    END
  END s1_wb_dat_i[15]
  PIN s1_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END s1_wb_dat_i[16]
  PIN s1_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 1196.000 332.030 1200.000 ;
    END
  END s1_wb_dat_i[17]
  PIN s1_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1101.640 400.000 1102.240 ;
    END
  END s1_wb_dat_i[18]
  PIN s1_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END s1_wb_dat_i[19]
  PIN s1_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END s1_wb_dat_i[1]
  PIN s1_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 761.640 400.000 762.240 ;
    END
  END s1_wb_dat_i[20]
  PIN s1_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1088.040 400.000 1088.640 ;
    END
  END s1_wb_dat_i[21]
  PIN s1_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END s1_wb_dat_i[22]
  PIN s1_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 907.840 400.000 908.440 ;
    END
  END s1_wb_dat_i[23]
  PIN s1_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 567.840 400.000 568.440 ;
    END
  END s1_wb_dat_i[24]
  PIN s1_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END s1_wb_dat_i[25]
  PIN s1_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1196.000 399.650 1200.000 ;
    END
  END s1_wb_dat_i[26]
  PIN s1_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END s1_wb_dat_i[27]
  PIN s1_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END s1_wb_dat_i[28]
  PIN s1_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END s1_wb_dat_i[29]
  PIN s1_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END s1_wb_dat_i[2]
  PIN s1_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 554.240 400.000 554.840 ;
    END
  END s1_wb_dat_i[30]
  PIN s1_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END s1_wb_dat_i[31]
  PIN s1_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 360.440 400.000 361.040 ;
    END
  END s1_wb_dat_i[3]
  PIN s1_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END s1_wb_dat_i[4]
  PIN s1_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END s1_wb_dat_i[5]
  PIN s1_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 666.440 400.000 667.040 ;
    END
  END s1_wb_dat_i[6]
  PIN s1_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 1196.000 344.910 1200.000 ;
    END
  END s1_wb_dat_i[7]
  PIN s1_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1030.240 400.000 1030.840 ;
    END
  END s1_wb_dat_i[8]
  PIN s1_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.040 400.000 374.640 ;
    END
  END s1_wb_dat_i[9]
  PIN s1_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END s1_wb_dat_o[0]
  PIN s1_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END s1_wb_dat_o[10]
  PIN s1_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END s1_wb_dat_o[11]
  PIN s1_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1054.040 400.000 1054.640 ;
    END
  END s1_wb_dat_o[12]
  PIN s1_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 1196.000 296.610 1200.000 ;
    END
  END s1_wb_dat_o[13]
  PIN s1_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 435.240 400.000 435.840 ;
    END
  END s1_wb_dat_o[14]
  PIN s1_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 1196.000 264.410 1200.000 ;
    END
  END s1_wb_dat_o[15]
  PIN s1_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END s1_wb_dat_o[16]
  PIN s1_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END s1_wb_dat_o[17]
  PIN s1_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.240 400.000 95.840 ;
    END
  END s1_wb_dat_o[18]
  PIN s1_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END s1_wb_dat_o[19]
  PIN s1_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 190.440 400.000 191.040 ;
    END
  END s1_wb_dat_o[1]
  PIN s1_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END s1_wb_dat_o[20]
  PIN s1_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END s1_wb_dat_o[21]
  PIN s1_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END s1_wb_dat_o[22]
  PIN s1_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END s1_wb_dat_o[23]
  PIN s1_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END s1_wb_dat_o[24]
  PIN s1_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END s1_wb_dat_o[25]
  PIN s1_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1196.000 80.870 1200.000 ;
    END
  END s1_wb_dat_o[26]
  PIN s1_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END s1_wb_dat_o[27]
  PIN s1_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END s1_wb_dat_o[28]
  PIN s1_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 1196.000 206.450 1200.000 ;
    END
  END s1_wb_dat_o[29]
  PIN s1_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 591.640 400.000 592.240 ;
    END
  END s1_wb_dat_o[2]
  PIN s1_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END s1_wb_dat_o[30]
  PIN s1_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 992.840 400.000 993.440 ;
    END
  END s1_wb_dat_o[31]
  PIN s1_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END s1_wb_dat_o[3]
  PIN s1_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END s1_wb_dat_o[4]
  PIN s1_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END s1_wb_dat_o[5]
  PIN s1_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 969.040 400.000 969.640 ;
    END
  END s1_wb_dat_o[6]
  PIN s1_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.840 400.000 58.440 ;
    END
  END s1_wb_dat_o[7]
  PIN s1_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1196.000 161.370 1200.000 ;
    END
  END s1_wb_dat_o[8]
  PIN s1_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1196.000 148.490 1200.000 ;
    END
  END s1_wb_dat_o[9]
  PIN s1_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END s1_wb_sel_o[0]
  PIN s1_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END s1_wb_sel_o[1]
  PIN s1_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END s1_wb_sel_o[2]
  PIN s1_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END s1_wb_sel_o[3]
  PIN s1_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END s1_wb_stb_o
  PIN s1_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 785.440 400.000 786.040 ;
    END
  END s1_wb_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 394.220 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 394.220 181.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 394.220 334.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 394.220 487.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 394.220 640.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 792.390 394.220 793.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 945.570 394.220 947.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1098.750 394.220 1100.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1188.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 394.220 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 394.220 257.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 394.220 411.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 394.220 564.220 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 715.800 394.220 717.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 868.980 394.220 870.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1022.160 394.220 1023.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1175.340 394.220 1176.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1188.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 1188.725 ;
      LAYER met1 ;
        RECT 0.070 9.900 399.670 1189.960 ;
      LAYER met2 ;
        RECT 0.650 1195.720 9.470 1196.530 ;
        RECT 10.310 1195.720 22.350 1196.530 ;
        RECT 23.190 1195.720 32.010 1196.530 ;
        RECT 32.850 1195.720 44.890 1196.530 ;
        RECT 45.730 1195.720 54.550 1196.530 ;
        RECT 55.390 1195.720 67.430 1196.530 ;
        RECT 68.270 1195.720 80.310 1196.530 ;
        RECT 81.150 1195.720 89.970 1196.530 ;
        RECT 90.810 1195.720 102.850 1196.530 ;
        RECT 103.690 1195.720 112.510 1196.530 ;
        RECT 113.350 1195.720 125.390 1196.530 ;
        RECT 126.230 1195.720 135.050 1196.530 ;
        RECT 135.890 1195.720 147.930 1196.530 ;
        RECT 148.770 1195.720 160.810 1196.530 ;
        RECT 161.650 1195.720 170.470 1196.530 ;
        RECT 171.310 1195.720 183.350 1196.530 ;
        RECT 184.190 1195.720 193.010 1196.530 ;
        RECT 193.850 1195.720 205.890 1196.530 ;
        RECT 206.730 1195.720 215.550 1196.530 ;
        RECT 216.390 1195.720 228.430 1196.530 ;
        RECT 229.270 1195.720 241.310 1196.530 ;
        RECT 242.150 1195.720 250.970 1196.530 ;
        RECT 251.810 1195.720 263.850 1196.530 ;
        RECT 264.690 1195.720 273.510 1196.530 ;
        RECT 274.350 1195.720 286.390 1196.530 ;
        RECT 287.230 1195.720 296.050 1196.530 ;
        RECT 296.890 1195.720 308.930 1196.530 ;
        RECT 309.770 1195.720 321.810 1196.530 ;
        RECT 322.650 1195.720 331.470 1196.530 ;
        RECT 332.310 1195.720 344.350 1196.530 ;
        RECT 345.190 1195.720 354.010 1196.530 ;
        RECT 354.850 1195.720 366.890 1196.530 ;
        RECT 367.730 1195.720 376.550 1196.530 ;
        RECT 377.390 1195.720 389.430 1196.530 ;
        RECT 390.270 1195.720 399.090 1196.530 ;
        RECT 0.100 4.280 399.640 1195.720 ;
        RECT 0.650 3.670 9.470 4.280 ;
        RECT 10.310 3.670 22.350 4.280 ;
        RECT 23.190 3.670 32.010 4.280 ;
        RECT 32.850 3.670 44.890 4.280 ;
        RECT 45.730 3.670 54.550 4.280 ;
        RECT 55.390 3.670 67.430 4.280 ;
        RECT 68.270 3.670 77.090 4.280 ;
        RECT 77.930 3.670 89.970 4.280 ;
        RECT 90.810 3.670 102.850 4.280 ;
        RECT 103.690 3.670 112.510 4.280 ;
        RECT 113.350 3.670 125.390 4.280 ;
        RECT 126.230 3.670 135.050 4.280 ;
        RECT 135.890 3.670 147.930 4.280 ;
        RECT 148.770 3.670 157.590 4.280 ;
        RECT 158.430 3.670 170.470 4.280 ;
        RECT 171.310 3.670 183.350 4.280 ;
        RECT 184.190 3.670 193.010 4.280 ;
        RECT 193.850 3.670 205.890 4.280 ;
        RECT 206.730 3.670 215.550 4.280 ;
        RECT 216.390 3.670 228.430 4.280 ;
        RECT 229.270 3.670 238.090 4.280 ;
        RECT 238.930 3.670 250.970 4.280 ;
        RECT 251.810 3.670 263.850 4.280 ;
        RECT 264.690 3.670 273.510 4.280 ;
        RECT 274.350 3.670 286.390 4.280 ;
        RECT 287.230 3.670 296.050 4.280 ;
        RECT 296.890 3.670 308.930 4.280 ;
        RECT 309.770 3.670 318.590 4.280 ;
        RECT 319.430 3.670 331.470 4.280 ;
        RECT 332.310 3.670 344.350 4.280 ;
        RECT 345.190 3.670 354.010 4.280 ;
        RECT 354.850 3.670 366.890 4.280 ;
        RECT 367.730 3.670 376.550 4.280 ;
        RECT 377.390 3.670 389.430 4.280 ;
        RECT 390.270 3.670 399.090 4.280 ;
      LAYER met3 ;
        RECT 4.000 1187.640 396.000 1188.805 ;
        RECT 4.400 1186.240 395.600 1187.640 ;
        RECT 4.000 1177.440 396.000 1186.240 ;
        RECT 4.400 1176.040 396.000 1177.440 ;
        RECT 4.000 1174.040 396.000 1176.040 ;
        RECT 4.000 1172.640 395.600 1174.040 ;
        RECT 4.000 1163.840 396.000 1172.640 ;
        RECT 4.400 1162.440 395.600 1163.840 ;
        RECT 4.000 1150.240 396.000 1162.440 ;
        RECT 4.400 1148.840 395.600 1150.240 ;
        RECT 4.000 1140.040 396.000 1148.840 ;
        RECT 4.400 1138.640 395.600 1140.040 ;
        RECT 4.000 1126.440 396.000 1138.640 ;
        RECT 4.400 1125.040 395.600 1126.440 ;
        RECT 4.000 1116.240 396.000 1125.040 ;
        RECT 4.400 1114.840 395.600 1116.240 ;
        RECT 4.000 1102.640 396.000 1114.840 ;
        RECT 4.400 1101.240 395.600 1102.640 ;
        RECT 4.000 1092.440 396.000 1101.240 ;
        RECT 4.400 1091.040 396.000 1092.440 ;
        RECT 4.000 1089.040 396.000 1091.040 ;
        RECT 4.000 1087.640 395.600 1089.040 ;
        RECT 4.000 1078.840 396.000 1087.640 ;
        RECT 4.400 1077.440 395.600 1078.840 ;
        RECT 4.000 1065.240 396.000 1077.440 ;
        RECT 4.400 1063.840 395.600 1065.240 ;
        RECT 4.000 1055.040 396.000 1063.840 ;
        RECT 4.400 1053.640 395.600 1055.040 ;
        RECT 4.000 1041.440 396.000 1053.640 ;
        RECT 4.400 1040.040 395.600 1041.440 ;
        RECT 4.000 1031.240 396.000 1040.040 ;
        RECT 4.400 1029.840 395.600 1031.240 ;
        RECT 4.000 1017.640 396.000 1029.840 ;
        RECT 4.400 1016.240 395.600 1017.640 ;
        RECT 4.000 1007.440 396.000 1016.240 ;
        RECT 4.400 1006.040 396.000 1007.440 ;
        RECT 4.000 1004.040 396.000 1006.040 ;
        RECT 4.000 1002.640 395.600 1004.040 ;
        RECT 4.000 993.840 396.000 1002.640 ;
        RECT 4.400 992.440 395.600 993.840 ;
        RECT 4.000 980.240 396.000 992.440 ;
        RECT 4.400 978.840 395.600 980.240 ;
        RECT 4.000 970.040 396.000 978.840 ;
        RECT 4.400 968.640 395.600 970.040 ;
        RECT 4.000 956.440 396.000 968.640 ;
        RECT 4.400 955.040 395.600 956.440 ;
        RECT 4.000 946.240 396.000 955.040 ;
        RECT 4.400 944.840 395.600 946.240 ;
        RECT 4.000 932.640 396.000 944.840 ;
        RECT 4.400 931.240 395.600 932.640 ;
        RECT 4.000 922.440 396.000 931.240 ;
        RECT 4.400 921.040 396.000 922.440 ;
        RECT 4.000 919.040 396.000 921.040 ;
        RECT 4.000 917.640 395.600 919.040 ;
        RECT 4.000 908.840 396.000 917.640 ;
        RECT 4.400 907.440 395.600 908.840 ;
        RECT 4.000 895.240 396.000 907.440 ;
        RECT 4.400 893.840 395.600 895.240 ;
        RECT 4.000 885.040 396.000 893.840 ;
        RECT 4.400 883.640 395.600 885.040 ;
        RECT 4.000 871.440 396.000 883.640 ;
        RECT 4.400 870.040 395.600 871.440 ;
        RECT 4.000 861.240 396.000 870.040 ;
        RECT 4.400 859.840 395.600 861.240 ;
        RECT 4.000 847.640 396.000 859.840 ;
        RECT 4.400 846.240 395.600 847.640 ;
        RECT 4.000 837.440 396.000 846.240 ;
        RECT 4.400 836.040 396.000 837.440 ;
        RECT 4.000 834.040 396.000 836.040 ;
        RECT 4.000 832.640 395.600 834.040 ;
        RECT 4.000 823.840 396.000 832.640 ;
        RECT 4.400 822.440 395.600 823.840 ;
        RECT 4.000 810.240 396.000 822.440 ;
        RECT 4.400 808.840 395.600 810.240 ;
        RECT 4.000 800.040 396.000 808.840 ;
        RECT 4.400 798.640 395.600 800.040 ;
        RECT 4.000 786.440 396.000 798.640 ;
        RECT 4.400 785.040 395.600 786.440 ;
        RECT 4.000 776.240 396.000 785.040 ;
        RECT 4.400 774.840 395.600 776.240 ;
        RECT 4.000 762.640 396.000 774.840 ;
        RECT 4.400 761.240 395.600 762.640 ;
        RECT 4.000 752.440 396.000 761.240 ;
        RECT 4.400 751.040 395.600 752.440 ;
        RECT 4.000 738.840 396.000 751.040 ;
        RECT 4.400 737.440 395.600 738.840 ;
        RECT 4.000 728.640 396.000 737.440 ;
        RECT 4.400 727.240 396.000 728.640 ;
        RECT 4.000 725.240 396.000 727.240 ;
        RECT 4.000 723.840 395.600 725.240 ;
        RECT 4.000 715.040 396.000 723.840 ;
        RECT 4.400 713.640 395.600 715.040 ;
        RECT 4.000 701.440 396.000 713.640 ;
        RECT 4.400 700.040 395.600 701.440 ;
        RECT 4.000 691.240 396.000 700.040 ;
        RECT 4.400 689.840 395.600 691.240 ;
        RECT 4.000 677.640 396.000 689.840 ;
        RECT 4.400 676.240 395.600 677.640 ;
        RECT 4.000 667.440 396.000 676.240 ;
        RECT 4.400 666.040 395.600 667.440 ;
        RECT 4.000 653.840 396.000 666.040 ;
        RECT 4.400 652.440 395.600 653.840 ;
        RECT 4.000 643.640 396.000 652.440 ;
        RECT 4.400 642.240 396.000 643.640 ;
        RECT 4.000 640.240 396.000 642.240 ;
        RECT 4.000 638.840 395.600 640.240 ;
        RECT 4.000 630.040 396.000 638.840 ;
        RECT 4.400 628.640 395.600 630.040 ;
        RECT 4.000 616.440 396.000 628.640 ;
        RECT 4.400 615.040 395.600 616.440 ;
        RECT 4.000 606.240 396.000 615.040 ;
        RECT 4.400 604.840 395.600 606.240 ;
        RECT 4.000 592.640 396.000 604.840 ;
        RECT 4.400 591.240 395.600 592.640 ;
        RECT 4.000 582.440 396.000 591.240 ;
        RECT 4.400 581.040 395.600 582.440 ;
        RECT 4.000 568.840 396.000 581.040 ;
        RECT 4.400 567.440 395.600 568.840 ;
        RECT 4.000 558.640 396.000 567.440 ;
        RECT 4.400 557.240 396.000 558.640 ;
        RECT 4.000 555.240 396.000 557.240 ;
        RECT 4.000 553.840 395.600 555.240 ;
        RECT 4.000 545.040 396.000 553.840 ;
        RECT 4.400 543.640 395.600 545.040 ;
        RECT 4.000 531.440 396.000 543.640 ;
        RECT 4.400 530.040 395.600 531.440 ;
        RECT 4.000 521.240 396.000 530.040 ;
        RECT 4.400 519.840 395.600 521.240 ;
        RECT 4.000 507.640 396.000 519.840 ;
        RECT 4.400 506.240 395.600 507.640 ;
        RECT 4.000 497.440 396.000 506.240 ;
        RECT 4.400 496.040 395.600 497.440 ;
        RECT 4.000 483.840 396.000 496.040 ;
        RECT 4.400 482.440 395.600 483.840 ;
        RECT 4.000 473.640 396.000 482.440 ;
        RECT 4.400 472.240 396.000 473.640 ;
        RECT 4.000 470.240 396.000 472.240 ;
        RECT 4.000 468.840 395.600 470.240 ;
        RECT 4.000 460.040 396.000 468.840 ;
        RECT 4.400 458.640 395.600 460.040 ;
        RECT 4.000 446.440 396.000 458.640 ;
        RECT 4.400 445.040 395.600 446.440 ;
        RECT 4.000 436.240 396.000 445.040 ;
        RECT 4.400 434.840 395.600 436.240 ;
        RECT 4.000 422.640 396.000 434.840 ;
        RECT 4.400 421.240 395.600 422.640 ;
        RECT 4.000 412.440 396.000 421.240 ;
        RECT 4.400 411.040 395.600 412.440 ;
        RECT 4.000 398.840 396.000 411.040 ;
        RECT 4.400 397.440 395.600 398.840 ;
        RECT 4.000 388.640 396.000 397.440 ;
        RECT 4.400 387.240 395.600 388.640 ;
        RECT 4.000 375.040 396.000 387.240 ;
        RECT 4.400 373.640 395.600 375.040 ;
        RECT 4.000 364.840 396.000 373.640 ;
        RECT 4.400 363.440 396.000 364.840 ;
        RECT 4.000 361.440 396.000 363.440 ;
        RECT 4.000 360.040 395.600 361.440 ;
        RECT 4.000 351.240 396.000 360.040 ;
        RECT 4.400 349.840 395.600 351.240 ;
        RECT 4.000 337.640 396.000 349.840 ;
        RECT 4.400 336.240 395.600 337.640 ;
        RECT 4.000 327.440 396.000 336.240 ;
        RECT 4.400 326.040 395.600 327.440 ;
        RECT 4.000 313.840 396.000 326.040 ;
        RECT 4.400 312.440 395.600 313.840 ;
        RECT 4.000 303.640 396.000 312.440 ;
        RECT 4.400 302.240 395.600 303.640 ;
        RECT 4.000 290.040 396.000 302.240 ;
        RECT 4.400 288.640 395.600 290.040 ;
        RECT 4.000 279.840 396.000 288.640 ;
        RECT 4.400 278.440 396.000 279.840 ;
        RECT 4.000 276.440 396.000 278.440 ;
        RECT 4.000 275.040 395.600 276.440 ;
        RECT 4.000 266.240 396.000 275.040 ;
        RECT 4.400 264.840 395.600 266.240 ;
        RECT 4.000 252.640 396.000 264.840 ;
        RECT 4.400 251.240 395.600 252.640 ;
        RECT 4.000 242.440 396.000 251.240 ;
        RECT 4.400 241.040 395.600 242.440 ;
        RECT 4.000 228.840 396.000 241.040 ;
        RECT 4.400 227.440 395.600 228.840 ;
        RECT 4.000 218.640 396.000 227.440 ;
        RECT 4.400 217.240 395.600 218.640 ;
        RECT 4.000 205.040 396.000 217.240 ;
        RECT 4.400 203.640 395.600 205.040 ;
        RECT 4.000 194.840 396.000 203.640 ;
        RECT 4.400 193.440 396.000 194.840 ;
        RECT 4.000 191.440 396.000 193.440 ;
        RECT 4.000 190.040 395.600 191.440 ;
        RECT 4.000 181.240 396.000 190.040 ;
        RECT 4.400 179.840 395.600 181.240 ;
        RECT 4.000 167.640 396.000 179.840 ;
        RECT 4.400 166.240 395.600 167.640 ;
        RECT 4.000 157.440 396.000 166.240 ;
        RECT 4.400 156.040 395.600 157.440 ;
        RECT 4.000 143.840 396.000 156.040 ;
        RECT 4.400 142.440 395.600 143.840 ;
        RECT 4.000 133.640 396.000 142.440 ;
        RECT 4.400 132.240 395.600 133.640 ;
        RECT 4.000 120.040 396.000 132.240 ;
        RECT 4.400 118.640 395.600 120.040 ;
        RECT 4.000 109.840 396.000 118.640 ;
        RECT 4.400 108.440 396.000 109.840 ;
        RECT 4.000 106.440 396.000 108.440 ;
        RECT 4.000 105.040 395.600 106.440 ;
        RECT 4.000 96.240 396.000 105.040 ;
        RECT 4.400 94.840 395.600 96.240 ;
        RECT 4.000 82.640 396.000 94.840 ;
        RECT 4.400 81.240 395.600 82.640 ;
        RECT 4.000 72.440 396.000 81.240 ;
        RECT 4.400 71.040 395.600 72.440 ;
        RECT 4.000 58.840 396.000 71.040 ;
        RECT 4.400 57.440 395.600 58.840 ;
        RECT 4.000 48.640 396.000 57.440 ;
        RECT 4.400 47.240 395.600 48.640 ;
        RECT 4.000 35.040 396.000 47.240 ;
        RECT 4.400 33.640 395.600 35.040 ;
        RECT 4.000 24.840 396.000 33.640 ;
        RECT 4.400 23.440 396.000 24.840 ;
        RECT 4.000 21.440 396.000 23.440 ;
        RECT 4.000 20.040 395.600 21.440 ;
        RECT 4.000 11.240 396.000 20.040 ;
        RECT 4.400 10.375 395.600 11.240 ;
      LAYER met4 ;
        RECT 145.655 30.775 174.240 1187.105 ;
        RECT 176.640 30.775 232.465 1187.105 ;
  END
END wb_interconnect
END LIBRARY

